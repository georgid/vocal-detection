BZh91AY&SY��(�s߀rqg����ߠ����a�O��������ݩ�z�P         �  @      �    ��Ӧ�圭 �        42 � �� iJ*� ���Ffyv]C��m�� �<     ��((
�8 �}�z� �iI(�Ȇk�6�V����Z*�9�aR��قڡiZ��= ��� �xm�]���C�����m��UJT��*5N�X��T���ڱ*ڬj��Qm�[[D����N<@Q'� >���V�6�v��SvУP��4-A�������)m@;h]�T���T�m�4]�K�p7�  Q� ݴ*�hr�*�[j�	4�uFE�BV���##Z4h���T�x �y�� e\#'kj�@���mD�lՕ[j�V�;��X6�ҭ�aQB���\ �w�  �M]jKP�ը��3�[%�SZ�`MPݎ��kU��MK�U�k6���x װ��l:�-�S��h��`�kWn�V�����W,DE�-�M�j��N��l.}<�  ��Y�j��6�D6�j�Zti*��5���j�mi���f��Իj��]��t�� 1���3��V�Mj���Z��[I�-��l�h��j-kT��n��J�.�� p  w�Ǌ��&��cJ�fԖՕT�SU��mQ���m�J6�vi�)q���&�        �CS� )IDF���@    )� ���2  	��  UT��7�5T�j46��ɣ@ � dhh��T	Jj� h  ���   ��R$%UFL � !�L&  � �Dd�i2OF�1'���m&��S'���O��{�{�?����᥹�KƸ��3���-�4~_�� � �� �� �QO�������pP 8v����������_�0���������������}׿l���s��9�g����(�����}�U�ӟ���" w���ϰ��D�>��n���zi?<�ϳO'D"��ݙ��9��?������s������y�?>��Ǿ���:�~u��r���QOM!"�g��׾]*�f��QF �C�?O�ӫd����z�>��3&���3���3���w���2�]��.�Pc����R���s9ˑ�۽���	���Ff'խ!��G͚t���Rm^������[
�1g�,s3�eK|��,��,��6���s��p��A���m���a��w��>�/HH,!s`�0DȊ�����\w��4�9N|�ɴ�ug�f�/���*T�g*�y�������WM����u.�J��� ����� �)ԡ$����E9U��>	�>�6s鮶����ׇiV7���U>��eP�˫	�Б�c��� آ�S˪6k� ī�rXa��	(E��MF��á"���t�f�l�s�8C��G^HG��a�2�߈�Q�)JR��;��)L����r_}�c����1�)�#<@�����L����n73�}�V� ��
�	/�!�*�
s,�<�����n���F�\�}���zx�x&f�{�/:Й����S���9Ѿ��J�ܥBR=��%�<-���-G~���N�.�W���^l��bh:P�~�3A��v<��l-K��g\�w�G^'�,H�T�'r�HE�m��N)�ޒy�Dl���<�O9:��LB�I�<�9��хq���t�Z�ֳ���{��v�N.u�hՒ�&C��pְ$�0L�-`t���Z�3Y0h�>���:�U�	0��������30L�a�睞p�ZsF�I���O�d�K,;���_0p�@#����5"^I�� 4�ik=���y�F^�����^g;�}�0nY %�V�A�ZB���=㉾==��Q��1�p����n�:uh�ټ��u7k�Z{���Vw�	�[a#y4�(�&��Wk\�9r]o|[�Y���7:(i��؝p�;=�ljo9,j�gA�������9)F:v�n�n���;7޳{�'�;��X�yy��L�K��sVm8ٽtM���.[��W�|ּk�S��������P` �� ! I��J�����G�(  � 랹����׊����֏ l�0�e��s�"J0h�Ǔ�� mrуA�ٴ �Kp�ǞTį_�<W�^��햬�w>\�G�R��՗�/z�B���� ��A��e ��� ��,���(�bTh�����)�+A�Ef�Z5��k�!׭k�fXW�`�φ:�?�h��-��`������k���9рD���V��~h�F�C^���@l��tlu�@v� ��E z,@���8 KeP�P��  ����v����mLu����ꃯU��`��A�!E W ��p�:��(�,���Q^=yN�z���c�Z��e�����y6�����~j��]W��l� $���]������׳���:�}h
�õk�P6%s9��hb�@�^���Ec��� ���.WR׏_�����
:랽��T�]�_\�1�;=���<�%�t��q��GX���U��z浾�&On��S]Q���ؓ�lۀ+�����z�ts��u���i�X6Zc��ƻ��t  �9��  � �[m
�MV: mZQ��e�\�U�`
e[�8W��o����^���e Ɓ��h�±:�=�>à�xt����0 �  � ��OL��:7*߀z�S�ۏG��#�hb��W�A�v��4 ڴ k� i�� 2��U2�  Z��T+h eZ  �n 
�� Z \�� -4 Ud�� V�� �h��@�ʴ fP\:�	�  r � `4B �p ( P0��Ȝ�rX��mZ��ٴ����6�UU���h��e�::�@s�jр6�
��hx�
�գA���4x]�� -r� �o���KCƽ�q��@ƌu��LuׯEu���t(�� 
q@ S�Q��	X�@�j�[hI@r`4W\�9=u�u���9]kx�c�!�ƃ�z�1U�c�䜒�\�ꃁÇ

8�rQ�PrcA�0I�I��  ��   �  !  @   �  !  �����ps�������F?=W?%����+c�b�^�|�W �V\xߗ�Q�Ӏ :,O��լQU��1�7jLh��5���;����D&�0������Eh=Uve�ȒtK@�[-  Z�4^�&ޏ���G��x�=sؕ�=l��r���^y���`���U�k�f| (7�0䕯{ܯ@w�*{����x�{�� -  *� 
�    �@ P >I�Nr�&eǯ�4�� �J= m���g��?
��z�úa�� �cAF�5�Ѡ�۹� w��޽x��5���h�=z����r�̥t��� �2�:��k��>r�/�쾊���jz�5�od�`�^�4 �� �U�ܠ���ܠ-�1�|�����(��݃��C��ѣ�P��_� ��h� �r� ����]��Cm�Z(��_��.��9<_��tz�)�ܡ��M�91�mV�: ��s �Pn�h( �{�p �u�_��Z���=z��x�Q�ƻ�{w�R�)R�)��`��`�ۃG��    @ -�P&{C�Q��l����@ 	��� �i���  p� P 0h��9�rV�P� ��8x�=������������ -���h 2��$�  Y�K@ �+(�e[�
U� �h ee ��@6�h 3���k�E6�� �� ��p< 3j� ��m� ��NPfU� =e��t ʴP�W PFZ S- h�h `Իk]�v� \�4���P�n��x��� D�    �  "  �    �  "  �   �k�x������ Q�? �x�cT�� ��  +:�_>k�W�c�<��р��(0k4x�� ���Ǫ�+z�~cF++�W�c����^
�M��. )��|���@UV]�rx5�:��� ����W9%�NP
��NH�l��u�����[��b���{�����Ƀ���汮|�G7�1���_=ϰ  ˹@`(�P K��j� o �/�� �� �Bեt��n�  e�( .e �$�'@a x*��֚*�Jĝx >�e�[ �6�P: �iÁB-��p
1O�����Fg��ڋz��7��	�˒���0w�E�uo� �,J����X:��}D��J!9�`(�׍��{u��/�k��������V�_
������~�0u��m�~d�TΩݘ��0y��7'�ߘ��Ǜ_,v�_L�uo��M;u�N����<x��{z�k�|��_Ǎz�Z�-~k��k3osuۘ��̺uL���Nۢ�����uF&ۍQ��[h�(���
�[�
��i� �k�s_��e�걢��5���6�=Pw0  ��  33  �� 30=(�ܳ���y�h����� nJ`�(�����~��]UWj��<o�� ~�  2Z  _ـ {�  �̘  ff  �� ;�  &�  U  ��]W�>k�πF{�<A�Tx �vU�<�����Q�y�%�� ��Z�4�̡���4rm�E i�2��e����Cm z:�y{��W�j�����''S�h��  �˙z�׃���ڠ�v�)����|���/+�xף�]��@�c�e���ǯ���{~�:<O3ǯ����������<�����ƫ�=��z 9�f�ׯ�X�^�Z  �֎I\�?jd~��'�hmz��1xR���4�Nr��}����y�~���	��~���[	�4/'���H�������z���z	$
~n���I�a�n��z���Sy�S�mz��e[2>lA�A�Z#�y���Չ��<�� ����@J��������C����	���Nyᾶwݭy�������~s�9���h2̶a���>N��z�ӭ&e�4��g�u6�ޞ�6ua�j�bgA���9�М��3X3�6v���h0ۼÇInq� � `�CR�n3 �RʺPFݯy��YO�u�/ Z{Ճ�ǳ�V�{��lo7;9p�1k�pgV���5��w��CQ�p�mޱ�N�ǳ�B��\j�w�]W���۳�s�j��TU�
S(ӟ+��i�Y��V���w���6nR��)J�ܥ%/~�9Yz�%��u�,��<�E�����m�.�B�Y��7������.a{G�(!��L� X�3�F�W&0X��Z� A��~>�(<��%ۚ�N��ﻬ�Bu9`fY��n���d1cD�3
�@@jfE9�!UQ썜8ܻ;g|�g��6s���~75�̉����I��G�8��Pqbg�ɔ<_�Q	 B�K����0{���+�j��>�Ͽ�������Y��<�}���^�k���Z���ڽ����z�7^��s���-̹{���i��m�ŝ�{")q�V���?�yo��9a�Cw�f̌��l�x�]\���7L��x����Yy��]����ɏ9�<���Wba������=��{�e�22e�22;������������FFFFFFFFFFO^K��ddddݒ7Y7d��FFFFFFFFFFFFW'r%W���q������������������ܝ�������f^/*��[###$��쑺ɻ$n�2223ݿ}�y������׷�ϵ���K���w���UVFG�%�Y��22q��2{}��ۊ�y�z�r�%�&��F�����#=/���ܝ��ݗ�F%仌����db_�.�#>���d���9/#"�]FC%�lmnG�^��9/#"�]FC%�lmo222+%�\s##/��ރjKUvm�aW��{�ow^`��כU����ݽ�]���yN�g��;2Q!��ۛݗ���ݩ�z�k�w��g5�r�����w�oek�n�o^kņ�޲+%�\s###~����}��=x���K�ddw'rn��n����22>���/z�ȼ��̼��M�O��1��ϣ&Vfc1�������������������vH�ݒ7Y�{����.2222222���3.�Z2>Ϸ3w^fNn����w��f�ּ�̜���#ҙ/#c������K�������M�#v�7g�{���������FFF\�����##"�^E�v2{�y9�ww=����������������͗�����������������������ɟVfc1���������������FFFFFFFFFM�#wvH�ddddd۪���Ua�^��u�fV3���^�Y7d���#u�����������FFFFFFY��-�� ���.�,[i�45���7;N�f��m�:��]��QY�w���X����v�7y�^��1���պ�&t׻���v�ovH�K�{����]}3���9����M���y$�ww`˻����K�����K��7wg�
p�@pPe�݁����ؗwv	ۻ�����O�N t�
��� �v����|��v� ��ɻ뻻���K���    	$�      ]�݀ 32@        ���         ̐         �� ���%�݂O{��.���.��I$�]��|��@}��]��=ww`�wv	wwa��D���zd�v	ww`�wv	ww`�ۻ�K̩��ww`�wvI$K�����N]݁.�����.�I0�>����e�݃/���Ӡ8(�fbK�������.������%�݂]��2���쓠8(��
p�@qNP n�e�2����wv	ww`�wv	wwi'�rH�}6I%�]��$�N t�
	'��aӠ9�> S�ww`�wv	ww`�w~�􍻻�m�݃n��w}�n��8ӡ������wv���m�wv	ww`�wv	ww`�wv=��)���@| =˻�S�:s�%�]��%�݂]��%�݂]��%�݂/�v>�N t�
��w$�:t�$�        fd� ���      32@    �wv     � 8       n��eV\���p��%�݃ns������.�����UQ���@| > S�:���.O�w�!���y�W��Y)���L;������so$�Gu-۾����a�{��H6�dΤ]��OX6�ib̰6��eZ��2tƯ�`��#3;.��3��hT�rd*�g[�l3]�9]�������ٹ9�gi̺���ڛJ��=�{gg]�h���q�1����h���{�����n���x��B�._d�Î�8�D�s�wio4�����h��k�%�s��v��Êj�9�;P1Wm\q�4A���z�uP��>N��1������剄���W<v��Y�^�b�xl�[�P�*���ua����m�S^G���9���jtF#���t|�v2%8��������Kwn�幪n�7m$����؈�ji��wh�Na�ׂ�]��mF���Z;��#2v4��ݼ��յ���;(��Yof�\ۭٻ���{�c�^�R������BD[ʉd���o72�n������Ӛ��wws���0�8�\�s1c��f:m�ͨ
�s�q%�Wh|*�)fv�t�;y*���~��J��~�g{ӵ+L����������^�v��������ǹ�s�J2���N��7�I��K��\Y�Y��r���޼�[���8üΘ%K:�ɘ�������o�9���ɮ�u�V��S� f^67B�7M�)u��gEZ/���fPx Y��&�w�5�dh5df�٪�F��Aޥ���m����k6��V���̖o3.Yoes��{]�u��1l&M�q��#�n�zfIIZ��ي ��Ov��°�F�@�ל�s�yzoOH�����A&e�so����j�YY.;���}���oe�Ơ�>9َ���n��7� [:��yċ��M�wX�r�����ab��ϧD'2�m�}{�vw�ْ�ܽ/F�\M������7,q�j|�âe��P���q�8·k�<��[���c�5�����ue��&��ˋR��=�����/�{2��\,�]�����z]�y����%��9Ǻ�ZՃ��٩��jC�u�#W�y�oaً�m�5�.�<�mܷx���Th1s$�У���q��{��h�ђ�G;�(��)ݞ����OWZ��-�n���L���+�
��\��+x%J۹/���Ll ��r��4��&t	m�J�/N��Z�x�8�N�G'��l�87����	�ۃR��ֻϸ���'Q.��v��R��٬Xrdv���%Á^rHL��;�t�O2�7�{χp9ݵr\9���m����_b]S��ɳ3Y�n�n�1[�uw$x���7h�v������#����cΒH�P�,�nd�f�R��XY����s�]��堬$��,qĊ�J���ÙJ�\�y�rP0,�-��0=ԛ��|*I����VӖ�Mdd���Rշ{>��JŃK�n���.Ү�.��޲�wD�L��H�wbgI�2�(M�]����Қ�V��m��tۊ��N�V���ZQ�Yv�=NӡًgPjw��9���M�=���17�{��q+%�ٖ(A�5�yZ([I%dn�j��^m���"I۬x�Y ��{v����N���9�`o,��cwfX������s0�<�n�n��3�,�ך�Ig<���2Gr�>xȷ��@$��B�ճ-�۰5٘�^f%5,�,T�]n������n�\Y�ZS7�k�ջz��u�WEHIg&,J�� �ѫ331�7lt�$���}���0��/�=��6����u�b���w�({1��w�SD�M�đ���� a@����w�5�<��^��7�d�s�jp�չ����m%4�7^���Ծէ��T�4��rE�����ͻ��dfeff22222�.�6o8��y�9��rW��W֯�9�<�6�`�ۺ������57Ͻ�o�E����������������������[{�tݿ#:���<�ַ|�n��]��݉)LA����>6��`ՙ��k$��&J��=�H���wU�m�K�ל�C�ܙw�*�x�I3nK�%K뻽����ꓯN�ٻ��Yw���5��J7���ڔ�Oj\��y��9�>�Y$� ����r^�׶��J���\���מ��ݭy�r��Wy�m�3ٽs��:��i%-���V�gd����wwrH�V���}�o�׺�����P��-�i�;+{R��m�{�5��\�bl�Sc�y�L��s�y�9���n������]�z���i%����ww����ܱ]M-�w��&�l���y����Ŋ�ݽŸ�q�oojI.���f�1�<ל�wn�M}ۯ[��7:�]�1�=�,h�U@\���[U�qwu���1$�Ǚ{K3/^f5���Ub�5�m��tq�k/[�Y��v�޼If�׊��o3s&���g'�4�x��Z�[W|�ݞU�'`4�+w�s�+w30^^^^f�\=�w�m��傀ud]4����o1�[�/p����9Z��ݫ쿬����n{jT1����X�������Pb[e>�7R��f$��Gջ83�/���Vŉs��t3RȺ�hM6����-$�ٰ�7{{4gR�uD�x��9�9�z�7�]j�Uڷy���{�ds6JX���z����y����V4Ә�ұw��[�;���4a��7w4$&�ُ���fg޼՝��U����K.�w��i�4e�텶c��һ����-�5E�7̒(�C5(M`;S%��n�s�}}����ʒ�2N��E�wn��y���|����)Ө���ɓ��J��f�]�m]�Wřh�=�����s�y���;,�,��N9�`�ݶ��n8 �$�g �d�+<�$������܆����}�..�{ϵ���9$��I��obWy�L�wZpph�I&�̻w����Y;&�ýw�D����Z�ͽ��Μ,d�N,ǐ"�g]�w�;¶�=�%��卜�t�W\���a��w��*��Ve]�}+35���[�bV���.���6�O��_#ȍv�̡�&�+7ߟx���"PY�Ǯ�)�p����,�'�5+%���U���w�ȇ�kl͚T\�4ۑ����u��w�M+��1�Mٯu�:KJF��;�2[�c��6��Q5[ط���ݻ�[�rq���_��dddddddd����V��+w۵�U{���y����{������|�ݲNk�yO5<��-����3k�yۯwu�&�_9�������&�gv�c'̌���s��VU��x�s7u�fn��wQk�a̻w��9���ٯu��s^����绻��9���<�	$s��ۻx�U�]����/qRQf ���O�+7}��Ƚ��֤�oey{�Ϗ�L$�xK�"�r֗L�-�ۄu���fU�b�m<V����Mmݻ�Wwn�޻U��޼��Ո�so^��p�'<�4��^��}��.�G���F�����4]ݱ|�s�y�8MٯU�w-�y��,�����U^F�{�UYUY�3����u������]�f��ת�*��3+]d���a(�"�!�����ڸ{��76-ۋYe"Q��7R�����������W%̢�y��]�>H���]�.��v�m)�~z�)�+��r�g�=~�օ��뿯���y��}�6�{��cI �X�̭��=d7	m����vfor�\���K9�w���P��~@�}��L}�[���v�� �UPt�y��UU@UU@ U@�$=��̻�ufEWn��K�����ς\�A1{�UR��
�T�\������  >�.}#7�mo��q��T͙ 9�۽����33J��=7ꪇϯ3�$�|sϻ�U� A���\�ݩ~��r{>��� ;޳=�{��U]��%S��v{�@���}Q�zK��~���N�7#v"-�f�m��o�]���+*��U@{�ӽ�f�{����U_O��;ހ _�330*��:;�������w��j��n䪁�O� �9ʨ���$����	=�67wy�[m��d�^�3`��d�*�����N���Wy�I���UPfd��e�A�S�:7Z�����FdK��[y���$�}r�޻�U��]@��&�ݼ��qP�α�݁�,ѽ:J��ۻ���ob΋�uT1ٌ�IlՋ��f�~ �z��>�̐
�v�����g=]�n���ɻY�f    �� {�{ڪ�ި����|9����\���U��}��o� ������_�H>!_Z���=�6$�q&��m$��ǢP-�]H�{�{���Tg�a�v6�=[���
w�Cj�]�w�j�Ya֖�1�6���q3*�j�{` ���|�t���%�q�K����ԩ�۽���붲�7[{�Y9��T��ɍ�C���IL���;;�wwy$h6C)�Mm��Ofg :�I'w+�rI�����r��IU@�����yΙ�$���k��qw$�_���]�9ό����  ���g�3����UW8���n�������� ����fmUO�g}�x }��{���o9 ���I*�d�綩 �UUUzd�   ]��&}'��g>��͕Q_UP ��ꪨ���wv��z�����|������  � s��9�=�'�$�W���� � UU$��� ��������T!5�����\������z���$�{�*���    s��6��w� 
��M�8�@w�\��UU9�������n�v��^�z;ޛ�wv>��%U]ԓy�'��T�C��3����-�V�Uv�@�[UbW xU{� >U�ހ�:}��}�B{��}�UU�Ip9��UU ���� :{�=�U�zh;ހ�{$  �    ����   ;ހ  
��39�p
������s�I����>��]t�ߞ����y���m�-Ks����b=���`�a�]�ږe���Za@6u�F�'�~�TD7�W����
�Oٿ6����q��������<`��� ���lG�}����?�?��~��~��~B���@�:����0�/b}��|�P���6q%Q�[����%6��8@��6;;Td�<����v
v+�4QElN�� OPb���!BR%;V �=���@|4��l�n��RA�0ңf�{CA�.�Sh�]�(����!D�DN�ঊG����d�9���x$+ў;K���:F3DJV�t��U%4�D��pA=�|�TN�UI�@�P�z;�&@ ;�	�B&��i`�
J �eY;-�A�E���0A��<�l.�9 �{H�
��0Q��N�1�G`� S8�/N���A�:v�f�4x��k�bkjV�ؠl؂t����3�Q�H�.��.���׹�hxh.�zGh�
�
�(�@��'���(b'�G��U�Hp��7���^���T��r�G����<�@�pUW�A<ª�I�1��:D{�J{DEGb�z�O@�!�)�a �dY	I@�%`(I�:I�!�U��7��=���{�0�8���Ik�@�%+�ц`��oi�Q��!�E�GzD���)!*R��>({� �&��(��)*���HE����@o�C�{en<X�@��B����(�G�5�����&�D�S�Ѓ��U�(�J��<T���@⽄&'��1v�z�K���u�E@P��W`,q$F�<WB%A�TE�(� B��C = `?��ߏ�@	�?^�6����j���z�hO�R�
�
j
h)�	JF�p8  �$!"$�ĥ)J��(J����(J��(	���( �(J��(J�(J $j JD "B��������)J���JX�����(JR�� �         �  �	�NBr!(J��*��(J�����(J���(J��(J��(�(J��(J��)
(R�  � �$ 8q Ü�  �  "  �   
�J*������)JRrBp�!�  �  � ��9!	8s��!�C���  �$!!8H9s�D    ���)JR&������   @ C�$IH�  D  ""    @   D    @ *�)J�JR��)JR��)��*�R��B��� ��Br����'!9    p  �$����9�Nrp    "    �������B�ZR��r  @ 8�)JR��(j�����  ��!9�N	Ȅ�(J��(J����(J��(J��"a)h 
 *��(
���RJ��_�吙%�4�P�%M
T�45	BR�ADU-"�%-JR4�%BP�%	BR�	I	HR��S����5���l]Vʫ�XlE�6��Q��UX�� V�
�3-�ZU�V۬�ڰs�U+��w����~�� fd�� �� I6p fd���̠�fn�>���d�˼��rz@q�����n��� v���UT��{}�����GP�M-��#i�J���K6i��ci\T�6˘�퐤 �.�2:J�u�ۚ�&-�fI]�]�X̎�v�P��ld�yv����v-n��*\�̂*h�7*����Ji�4�ٱnQ�]�ې�^:��ŋ46�0�P���b�n�Q��[���bc!38�]۔��֛[��u�+4�Z�\�C"�!��AG��=�iPW�piݍ=ȚM�j�l�\�. C9��#��!!)6XIl6�s778Mʸ�3�����Q9���覜GB*X}#�h��[�뺕8�[ݚ������I�8큄�g��e���Մ�Q�Ӂ'$HѦMh��ιG��ݳ�e���"5���Un����G�[ >
v��)�@WN� eO>�CblA@�qO@�G}�4�U*iD�p_9�|�u�(�C	�C�H{��]D�|fO�����lE��q1q�Q-��<�ꑈM̆�4`��S��ux�%��ȧ�B�t�)~D:@E�9��̬֠�f�Y��\���A\�@O����s���y��������{�~�[ᆣ]a�h챰(,`5秢I�.��w߽��A��Gid����#l8t'����eh�pHLt��Fޓ��bBI%��1�c�0�,��0�~z^�v'�z�xx>�LbDi��#v��\�NN��9$0������C;9���ٽ��$�w�씐�۱�q�H�-	�S$
GA����a/#����f�����Fpt&�"a�b����E���A�kM�A�&M[���611�.&3/;�|�MTFh3M�}�����œI��K�m��7,N�ﾞ���=6x'�.�Ii	14�`���qq7Ώ=���8}}D$�O@�o�w���@")������"W�7w}��cԳG���q!�$dY	P�1aXd$a��B��.G�P�Ŋ��thѾѾ��7λ<��}����%�4�l%Ą�Y��
�����&0� �j���bǰ�їM�"(�VXР*�1�쭕~3D������,o0��B<=Ŝ(��Y�`1�����ӽ���S�w(� }wsi)z�Kͻ� rH.�Y�20(JG@Q U��a2@9Ntu�jM'�(zN����}�x�<��@{SD�=1��F��T�.P��{������)�Aw�f�N����=#^�vFzo������4 ,X��}�0`�D-�Q�!�ܗ8��������(x��OBHB�I�.$�!�<�sF�9�F:s|��k^Io��zD�"
������������������z�_�� @0��uT�n�бi�����>"H$i`5��< z"�ïb��@�>Z���M߄�g�,I�H$�"%�5�8톉wI�'ҩ�-�kVά��3\��Qk �5�X��T�Pt���׽pp`�;��vj��)[�O4ҁ��0N01�t|�?YTbM&�2��[e+�+��~���{�:�?_nT��m�.�L�i�@�B�!�m�����傭'���$l��׉��q�:�0v�4���.��N��,}���{B�)UJQ��B �@IS9�]s35�W�wo33̍P�3�5ƪ��kLʺ���}NK�*Z��ʼ0A���v6���k@�M��7D�cOכ����ݹ�1��pVwN�l��ꔜ�R7Gj�&N��XeIcPيӻ��Ue̝��6l,2�Ώ~���:ﮋM�M~4�u�\\ۊ�^aCޏ~=�}:��}R�BE��F�"Z�M����%��
�7/0hn�D1��K(�K�*'�(3��*蓨����:������;B�z�L��-�x0n��%��*��ɆkcN�	xx =�*,^�ތ���v]۪���SwW���cv�����<mM��fȳ�ݺ��qV���F����~�������o���^lg/+j�r�sI�4��"������wpT��u�~(ԔHT�rB0���Y�������W������`��};��Au?��'�(��D	T�*i���s�ݒ���R};�n�u�+������lI�u����޹�fS�
��n�d7�6j�v
j)l���%\fν�V�{�{s7}��E.�Q��c���TD�r�S=v/6\L*���VlM���I�yy$���N����Jm1���% UU��O|��:�~��6�c���������f\Mt(�땵�b����"ZMy�(�SP��x�ֺ�f��qu�/mL�*�t.�ņ#Y����:�h�f>����kE�5�"�(�P5,J���j�L��HR�r��F�ys�n����}���3f����| ˬ�"�b9򔖋�_�A2[�UF��Ye�v��͘B�uw�v~��>�M-��)��L��F�k�r���\���x0t5y�¶���Mh�� �+��S�e�v��aCȭ��VƑ�A�c!/)x��t��\�P���-�\�=��˽+��U��F�j����,����F�`�zش�o)6[j;g�moI����VC�3c�M�]P�~��)m��t%�ٝz���؟BM~�v����"�m��q���)���F\kSqฤj��f\���iqZ��y|���f������-��:d�U ĈJ��9�Q>g7��45*�J}{y���H��5��%��$1T�{����ٓs;���F�aʇ�
)=��4w�"��4���!]��#�� p뗒�p?h�Cu)����-(s^e��ĝv�p@n�4C�y�0�T�[OfR�%X��o��]R���5W#j������/,��f����3Y��f�ؠz���}�����tte�pE뱱p*��7:��!4��lU�L��j[�ܷ�nB�rs	6(��jg"�j`b�C�HŘ0�N��F0��w�fs~w���Z�̧�`{ufmr,fu�K�ٳ�  =�y9�*����NH�x���y�q�R�*r�+���ؕ����m�n���[ǡ�ױ�٬Q)�l������nw<���z�w^ԩ�\�"���KN�H��U=�ޟh�B]$l�b�TpXR���.�t�����{�T�l;P��P_�9�U�*�(�dPJ��6Rim6I��
r�i�*%��B�^�[�J8,fA�%��gY��[ۚ��GJ��͑G�{bde+��
)%AP��7B&�\��5��>r��+̮�M���Y1���7�s��z�ܭ��[yR��՛�B��B�^�S�^��{ε�n/��X���ӷ�ۊm��F��+J�"�}��2HzM?^p�˒$� ��%���U���e��ʧW��Ȗ����6Kl(.!�nmn��-[,<���n_����-���P숂��	(�$Y��&���͡s�� ���*��ʹwX5�WB�$�۔'wX��*����j�^�tL+Ҥ��Y#e�%��.�V���suH�%�{������=\���7J)����V�����קn��Ӡ=N{�~}�k���cv�\�Uw4)��2ԍ���&��Ǝ��ܰ��SU��]r�e���h�n�*-Y���IZ�s���cm�j2��ɦ�H^��l�Rq�.��Q)�b��@�;\85�v�4}����K�Л���K�l��!�n��K՛Bg؃K`����a Jad��l��ݼ��gDVm�+�v��ۊ�tcGY�V {I4]���I[�����[�ܨ�k��Ƿ�N SAXEՔ�@TkG׽rC�0ݩ��G�q�]�g;���0�cn�ת��y��=��l�۵���{�u��y���\dPp�i(-�o�Oz�{֗��״��==B�5b���.�E���c(`׵>�iC�����qg9ȴ!�P�G�Bْ���fc��U����h����7�tiA!t$.��*�d9�&е5PKvtL��ߺ<��M�Ώϗ��:��&׿Z.���5ڎ���}Y���������[�U��F�Z���J+&
]��{�nl�������n��N�ة����V���4�lD1�b�������_t�Գ���IZ����D��R��_���]��[)ے)�d����՛1{ywxn��GK��v."��-�b�p��"�[�b��n��l6�n����ܫȩ����x�(�=GJn�GH�iP�J��L��������w�@(E��+��O{y�$|����)(����z01����,��Eݻwٵ���;��ޢƮ9;���%��l�όwV�ƶ]:):ݼ����I�1��id�:��E�ͫ�'&�HR�w��D�������1�pF�l���xgY����o:
�6�шXj��_[��DՅڕ٫�-�*$�8m{�
j'6����zQ�cN2Ra ����!I�@a�l쉰]���g�Zp�Ѐݽzr�!�\�I��U��"�
Qk�1�;w�+�VTaE�emY��8xZ����t(I�.j�*$9����W[�<?�_��p*0$����#)α0�~�j|��18�:sA�j��N���<�\�!�HH���b��SN�O,8��a0�����4�BNR1Ѩ4�ƍ�hBp��N֝�ٻ�R���X���4�,(��H���A:����i'P�K�q(lh,pc	�iq�ɷ���UUP�h޶m:%9(�»Ղ�T#���*�V�5�����S*����p�UUUUB�l��/C��Hp J����FN,8���=rK6�8[,�8ɑv@$�0�[��CLS_]�n��2e��/UVض^[e�-��.\�rX�����SH�Be����X�I�Yb�J�y9��8������K�z��a�;�R5C�P�Rѐ�^l�[q�$��c�1/.Y7��F��4��Aa��9fI,�,M�j��A�oP��;��u��k�u?���e�ʋ���GÜ�9��9�l�9ͱ��6дL�Fm���K��˜暫u�s���v�9�r���0L�M��\� ts�� Ύ�f]Cs��sa�ҹ)�t���s�����wwrg{!N�e���$� \� I#wf��3�$�f�� zH�$�y���I�U��I&˻�>� {�@�z J�-���\�V`���i�r电���t%�(&�j�1�6:]q����Z�[`"bź��h�P��L(���5MF�ile���2��1���%�W��l�:۩M�ʄ�����)M ֈ��8ЦY�қZ�5n�J�a��6�6���쫶��+Z��� �!���]K ����M���%(�K�R�aI����Z��h�\W���uΆԘ\%���:Vf�b7R:�h��̢Y&ŮV2�7Ja��iQ�cMq+���]\P�t��%sl�_�u��Sif���i	e��m�p�UHU�i�B�KF��B�!2�Q#bg"��d��,؅�1���GM�����4���}��}g5b/w�i�[-���kb�+uoq��/3��Wz�w~�������hd3�ZVU��;�'w����6��Z�DS�)l��s{�[2 �+0�m�K[j���Y��<�I���7����wn�7	���l�wwg
�����=I�IfdMM擖��㈆��Ր�	'��Cb��!�]*:�t��	| ^"�x �L0�$RQ|TS��LM"|U4
�>	��� �*�ӽ���k�6��i��r�/��Яe<�z�}��nxY ~   ,1�����͂_I�nI���O��"x��J��:|�L��f'�Y�:�p(:�����9u9�s@�0��)u&���G%��9�>u�˴�;�	#�
>����Y�Dz�� �I��;��a2��[4�'�a��W��;������k��F���V��{��Ty7 	@�O���7p�Z��p|��c�9O�u�3^�/GX7Yb��J�m2�u';��>O�nN|�䛏��Z��>O�9��J��2���uET������4��Y�N���}��h����Nj<iJ�TԁDI"O���Й Z�~w����\�`��7]Br2p|�j��3ʞ�ԟ<ǫS�{�����oG9\˟$�u�l�F��t&F@�j��~G��;�	�&̹��kW�~s�xr^�`�:�W$j��:�=��`قy��ϑ���z���uf��]ϒ=��׳��J1@��@������>�q�!E|��מ�͇r!$>3�s�����Y�Q��6
�řK!�[�����$���;Z������fRfU��
GK��"�[�k�kiH��(4YT#��fm�_�W��Z�e��Y��.�5Q2Z�W+��o��A]����c�$y�{�ed��}�=��i���E���Ƅ+�LB��g�0�{�MOq���Ju�Q�O�$��0	R�86�%�#��Mu�v��޵�ߞ�Ҵ&;����r<����%;#�ܚ�癘f��Y��
$�  "�
-;��՚8z����:���>g=��$�\��s;�N>�$D	X��qN�"�p$���G��{���A;C�"��Gʦ�f��F�((2{�|Ǩ��f���	�!�������إ�>y�S���A�>|��qDx4��[>wDt���vfuk����#Ws�&Bu{���/k������ T��ٛ���$T*{�9݊W�N�@|��Ǳԛ���qlXq>L��\H�&O����R����I���U'��y��&���	����=G����}� �WP�P,���>ۺ�T��L�s�G��7'���|��>K��E@ﾻ�R6��ݖw�\��p�6�u�R쯾_%>dq�<@����(ꞥ�;�,���9�Ϝ�f��gw��s����XCL袚���C�t��۪���{.%�+Rd�G�G3,X�a�k�FA�t�q�`2��٬�w���/[�1�N�������
i��!),(�m��7.�LD<H��wF��p�!�s�jM�Z��%��9�{�]�H�|(�OE�<�
��ָ�]u�Y������!�%3�Z��^��wo��|}����� H$�O��~g͇r%({����]C���7=�#�=�R�3A~���i5<�{����
>I�}�:�b��\�3�j�_#ϙ�|�����I�>�QG���dY�9lܚ�Ro[뮺�$�+_=�|��u'R��9�Q��x��Y��z��i��o:�i��"Ϥ��A&��'�2w�f�<�s��������>Gp�DH�=��M�"VbX�ZQ4\y
A,����zxJ֢��O�Ro�Ow :�"��{>���f�;4������ݒ6AﳧWm�Y�n7������#��C%<���!��ޱ�Q��5'\�j�`��"xǺ]_f` �G���������Q�dz�kA�N'�8�	�R<(�Q� i���@dT�U1�%�w]��0�7+ͣ."�ݬ�N�2G���u���&2O'[�5ܛ�S�&I����=.�h(lݛ���(��ߟN��N��uֳ3�}�P���o��ԥU��|������i�W�̍4G�佻�@:�2Ρ:������V���xZ�2EEE�>���NMfk��F�m�#��&Lu��/m�Dk�B��tt��`�G�,��%ԽW�# r����-/sͼ�HW"�k�CM,�\8.
no���>�y#n���V;���/�^�X=��FcBe�jy�\j��¦q��mF�!�l�W@��g6.���62�h���QI����xM�/x�W�r�e�4�7>ېH�TfF-�1�������+���t�NK$7DP�?n��j�
����k����AىEDX2!"M҄����z�����V��d7����×w��s3�]���^�x  <���8i���B�b�6L�P/utBTUzJ����������9:�+�0�:)T�#�tT�� ~_�~��P�Y������J �"U�������V��`�
5�F�"�J(�l��\0��?u�߿u���ޚ���Z)(�b^�P��)I1���tK���_wf]����z��G���_�ՓL�.�2�ڷHOZ,�#P��P�3(��TY�;z���m��Dh�)��*���(�,��U}��y[^��ػ�ܩ`͙���0�o�Q'f94��񡻳�(@ �n���t+���WJ"�RW;�S&^n���R����ч
��:ӵy{Or챊�xˁ�r� �ʠ��=s-{��J%V���<.��?��k�Hb�.������؅YXkp�AR;5�E�5ͣ?����{cZf���7�Knڎ5�ƻ�1��A7�~��o���4��6j5�4I������-
��Į�&��,��*�т�%�}+�jՔ �i٧U�B�-�V],Ĉ'�~��5]�.'bdZ�cmGd�G��?w����\YL%M/�]o��Ո ��Ǻ*i�Fإ�F�+�����]P֪��Q�����R�!�e�v�ś(��*�]���M�+0ڸhV�O��5h�x�η�ze�`�t̨��.���5��s�)vdt��=�������i�X� �m�c��CnŻ7�n_��ͮ�jP�S =B����sfo�C�0(!��+�W.m�WM��x׷؝G�_,M{mBa�ic(�
%��O^~;�Lf��2�bP#D
Α��C{�Ej�;���vn�ML�s�&՗S�)f�t՚�r�'H�A$5 Ioe��$�u�u�8�eՀ�� �)�(��E�VfM�Y��gN�w`=�]��UUo��t�$��e�i0X���Vb�{=��4`�S_� N���>���BI���@�l����ݵ�ԦD�C�׉҆{��IT=��$P�ov:�80/ nu���GT!w7Y՝������r8.��u�L�P�4�͑�-E#KȮ�c���x{���\��|�8�]�����mnDm��f�"�{�xx
Q�ɦ"5�-��/q\���������ؑ�mw����fB�y�DVYu1t��'{[�.
w����)���q�=᧺RTdl�����WZ��_ Yl�p �[!٠(
��2�7��՗�1��q�������t���75׀:\��H=�Q�ت�2��DLױ�Gx )�n�&=���Y��?cu�P��U�OV����<=��u�y{���������"�Є"ᷛ>����t*fR�lq7Q��=��J"�a)�xz[�|��9�<.;����G���UK8���˞��>���>��,PI_G ���y��@!^��C�{��G��um�f���m�XWFU쎌;?)�i_ۿ/�yXb�3��ΣmۭT�3ͨO�{���#��DǷc��c	�g�hڥ[6��Js�NU�(�iɀ%�[U~�[Í��#�QK���qF�k�	�W'w���=���}�P�
CH�Yu8%s	�%�*ϯ���x s����#!�1�|�7?��@�ÿt�:�7��Y�ۈt%EW��4�e�؂.'���EE�S,`_	з�v��v"j��㜻Wu+q+{�*T�n����x{�1���h4t.=�EZ5��_Z��ڣɕ(DX�J�j�˒��'<y�TH��jl�_U���%W��۫^T����WHnX��'w�(H'~xx]U�-�|�IE!�tFM�V�#���s����>��ɦF�Xv�����լ�S��W��#�tyP?yגI��w7�����\��}r���J�"a�^��@к���j����7%�6u����T0�n�k��v��|p��к'�Ѵ*��{Y���ɌQl�((*"dȫ�b.0�M� ��|{�.�ޯaf�67qV���­�j��7x�E�LWQ�;��*��O����lY�v��;�:�p�^��!$e��B���\F�Z��ZJ�L(:˼�ַoZ�0ѭ�
]�hl�Ur^ �+�v�;�RI+�~Ǘ���I!�\@#]ۥ�]��bc��l�۱K5��]�X�*�,�D��%�R7C;j�I[N�a���>Ώ8CI^C���fe1v����Mj�F��t�UK\K�A�٦#�:6W�F�2˺�lu[l"�䵇+T;��!�bWk��ɁP#N�=bE��d#�BD���6`��l��5}����a�+WkE���"��\�8��-n��� �(1'��1zx�Hp�b�-Q��ʜ��� ~��"?���å�
`�J:إ3�C��x{�jow���S��� ������!0�^ėԄNu��
������媊^��p�m�l�*_{�|��� =��,�[b�3	��LTꉀFE�O�=�� {�f��HQ��|m%T(ɨSg&�T�c('�xxz�����>����vk��W6jmB4S'��x{��=����O}t �^��*�1{i0܉� ]�0�� �0�#�I�6a���O\��X�����g8�ݘ�������}���ΰ:��)5P8d��9�vF�s����YbJ!e����L��G#���{8D��
$�z�9�&��$�  ���uޟ9�w̼��Z)��s]j&���P��10�ɳ��"x@�T�99T*h�69eYR�UP�@	UT�{!�@��4�*���DթE�����ʄZJ�M"(a�6�T�A���*�r  s� B��*ʅN��n���rH��HYP�����}y�G]@���"#�U�R
Ѳ���7���d�r'0NI�: P N   9�1��9�uP� �����a���a)���EMA�����6vM%wS�UUT(�wҤ�,��~q��;�GjM�fv���˳��2L�3�1	;+���Y*�r35jN]]�<�m�<L�)#3��U���)��՛*�:;����s����FK%�\���m��!b�a��*��UrslFՊ���m��\���t���=Y�Mu�*�V�����AY�7G�� ��: �� �$���e�����ْ��)�߻�����$�>�� f�v �� 6��U`���o9!:z����uZ�K�;����v��ف��%KAIyI���Sdt�j<�gZ��M.RT&Q�i�7)�����ڣ�6�Mm�y�e-#�Z�m�1K"��6�嵺Գ5�^W����+e�"9pX9BkY����bmQղ��V�Ӻ�ً͒�9��wfm/�m5�e�n�R�Xc+VYt�:��ep�,�����★AgEw�2�&fK��'�`:l"�e�5�є�=�]��-�I$Z�)��;���Ss�����H��g[wzOXxz�$ؑ>��ٶ:�>}Av���ݢz�6�Q��v`#	���������G�H�C(�D�T ���W���ǻ7��Pv�$�m�ݷp�4'E��l|&��x{�;�{ ���D�р��#���H�E��6�":P���O!D��  ;��̧�a-��-�j��&7;�.K'-�הW�Y��.Ye�a�jLJ�
��`)��\�����d/�3+37��"�T�����ӆ~� =�����a�zM���<�a��Q��Z��j(}�M�xp@u�}3�ך0���>���803#�T������b7��z�*_��.?��UKغ8-R�޺�{��<Tq�f���&$�ȷ�Z��Y���a�	E�g.�b�$f�
g���`�#,Td]�����΍�B�r���E�;�A���Lã��!^fW����҄"�e)�l;BA�u����P(������=i���C����ƫQ��>5j���de�t�N��q�H�\��r��������s�;-�ƈ����[� ��[�[��Ao����n��MC��3jgI%W�tT�2:D0�+��i��TP�F;�D/-@khn��V��M�q]2kY����νC��l�0�����	kkpzp�]H���NHE�	�j����t����`�G��hSO�@D������@4 �|#�RL��D;�]�˫��ؘ,�^��RI�$c�UU��v�w>����$}L��C�3�P#`���ċ��߯��큲��U蘀嘥o`9��1��	+��/'���`T̊�H��*�yI�d&[*D�X�������4�ɴ \��@�00�����;w>=�}�xi�8��!ӫ��Sq��Z6e�~}�+	�d���Bk5ؔ6�q�b4�}w=� �yLL�Z��}��B9��}�;�v���Mc��}����H��=�p�D]^����:��bcq�_џ�  �����}� G� ��{ߕ�R�]"�߾q���X4�+�� ��<Ĥ���P <��� _\!eL�G@�z$�J=n>�[w~�/}���ʔ��Y��ܟ@�ݑRLh��o���l6�b�\�74�78���b.m�������A�KP"� "�HP��*D��
���:���Ӟ�"Tυ0I=�%b��تp������7�����/��	���b�̂~10�ԅD�� ���Ͻ^>���,(�W�=B����7�;�M2~����
�R��Q�Z��I�2H[��a_���������$�SI������L>�k2x�En��f�`$��Z�q�� i>����W���p)i�-r�J���l̝;����$|n�R�L�W�	
��+U��'飗;~�H��/jFm"c׺��������o{@��J���f�h�K��q�8-R�O	XM�+������g>����B�=�s �#�"�SR*�K�	�N����6~?��"!l1Q��6g�*���iN�l�Z�X諲��J C{��aoJI��8N^�i� �bR���u���(i�Vl���F�L������z%6��N��[c*k�<m̦�ct�0ML6֍`SA�S+�߻�{��P��Q*�m�9�$�h ������΋�#�z��ɚa�*��E�0��bo��ê	�M�z��u�I�����A�D4㾟���ÊIf@"�X���k�jo��s����D$�A���B[P�jUz���=3���N�t�vh��G��i������	$�Cb�!�b7CJ�2Q��U@�`f����;3����ܧ����T`B�E�7��}H:t�h��X��m��I�&� nu& �%2V�=��3)L*	���dAg{�M��Dʚ�{Y��������D���Ũ$�|����t Ù�ޣ��X6�1y�0ԉ�$�i:�X艳�a�^5캺k�L;��%���^�W������~�J�kp��c�'A�YJ�-�����]�Iɮ��'f�"ڤ-�B��GGߏ�u�v��W���]v�	�P�[4`�s�.sxة�`��kLlS\���R��}�~��ޟw���_��!/R��!�BpX>W�ݝ�[�P"͠��b�$�E�n]ED�q�]��Fܡ�(�\�}�n�[Bv�̺A���sFf�� ����#�J�@�7�E�m9�V1��;�+�j�ٌyΈ�<-��U!ڙ��۝�}�w��x1p,]H`�T"綥���m	�%��KAgoH�����}�05��0 �*7�S��L� <	��1���k�Bv)�#M��Y��z�P�a
AR���YUtY7��!목�Gߏ��i���|
�^�Ds:���W��A_�����G 9��
&�w�=w��Hq��ݝJD�&%jⶓ����=0hV�/ά�B��{k���	�6�����W����fY%j��ݻ��ЅL��ݒ\F�꺻j�� 	��js:	/eC�}p7�EH�A#��T����ӷ����3�=�3!�Yp�@�W2��[6��׽BA� �_�=�"��7��洝U��R��]̥7v,)d�i�M����cI��q��r	���ŨS������Wj��F��A�-���i�.�P�c�ʶZ�B��S(�L�n7]m��[���b����ߧ9�'��2ū�ٌ�B�r�"�Z�{����sY�N��w@�0�U륏����Ei�Φ2�����i��:��׷������V�ўܷ�Da���U���x{��{��������щ�|��R�t���W��&�R�R�rS4�
T��	�z��@�����������ovU&n������f�T�&��ų�</��x{� d���Z�U�uD��esC=��tp�" }��wG��{�1�ѻ�L�#���1�D��P�l(��7ۢ�&�tBl�L
����f���Z|�\���!��t�h!qWq���Ʉ:����h��m�t`H�y*�ف�Pו��,����,~_}���������#.m�7�Nn����A��Ց��M;�������؍݈�-Ӥ���i�!���xO�UC���"(�l����"�*�Z���cnW� T�����{� ����C�
��M2d2p�ꚀA��r7k�2fzX��s�r-@��!tUy83I�H�^P��t���1\��ȕ3 ���X�"�|f!��!�($�~����
�yvpl��� ��W�ڛ��JKbF�u�6<T S(*&m#bK*�,����rZKj�%6`�.�֐�vl�9��Ѹ62�e��&�i���ڕ���+�ݝ�����g�m��P��AyM�� <������: +�3m0s��e%)��*�Uȿz��]>�y澚��Ι�/K��hFk�2ZQ���#�b�A�����IG���������읇N��ֽv�����N�Ȏp*�t�'LLz�%�0�҂wV���C�D�fL��h�Y�.lTZ2@��}�gW� {�T��vm�Dl�ɋB&�jP# ������� ۞�W�_A[���Zm��C/���4!�Ru�\���6��z��=.�	�\g��xq��Ԩ`���z������xxQ�r�`@<v�GH��^!�hdE̝~Ϫ��K
�Q�Kl�/n[&T��tp_��&�PF�V��LT�MJ�(2Zg�����j��:���-C����ť������|��A��FHd������K �f���
�Ɗ)3��~:�'[�'�}��y�u�m���ι�8eҐ2�,kr�:l�0�w�}��ߏ�x�;w�W�������L����l����<�	Gv:�� ���l#�K�gws�h��u��`��<�H��QL��y"��L}��n�ux�|UY�CB��S����?vOϬ�ޒ���T�ڠSr�DĝYj��ϐ�"<�ъ�����.������j��6���[�v�)R�ۗ������� �10/�K�a�a
X�{�	�7^�|�&h��q� �u񻨊G�Ma?~���DRR��A���X�SSksQLk������{n��/��P��]W�=����*]�Ǚk�Mn�j�&���$��Փ��#ᷥ��� WT�2>PI퉆��Ӛ�m̵B���^�l�������%_��̹���u�!X�f��`��)!9�i%��@@����|+c+�!RIg]ݼ��25��`��ݝ5J�4z< �Us��{�Q�Ο���C�Y��둑bz���޽����ݠ����Sp�]����Jud�G׳��b�� ��B�&Ó�еtU�i�؝3/.ܩ�H�Ϻ@���=��*��i��A�K��_b��P#�}��}�捕���^.�Ʈ�!����+Nx�׆&��׾�1v?1�,�ҵ�ޡ�E���8	}��ߠ}�ߐ�� ���!��Q��'�}j�m� �S2�
8�"XQP{;��^p�1GtS�)���h���"�on�o^ <����R��#���)bh�A�����K۾����O�r��VMB0����Ƚ-���^V���a��t�9)3XOٛo��t�&4�]���X��T��ֵ�bf��5�-&o[<��΋��,�ә�/fo4S�:8�R�)8�3N�l̔�c��Al5�R��5��V0 �
�.�	��{I!���	
&!�1��(���jQs4��wѭ- �bq �o��,���L~k��Yk7�j�(��S9�s�k�[�s��vÛ[\������L�ΛFXlջ93������l��r�m�s������9���9�d��E�s��s2Z�R���\�
#�������ot�ӭ��l7�Y�2�$ I �@I��30�����̐ {�@s����b䐓;�� >}'��d�I �$UU���	���}�j�UUՓ%U�LB������W6k�M�8�J�IClnU���n`ɫ]�͔�H���:���6���[4Z�۱ (���b���	��CY�i�it������`�T*��X���3���x)(�`%)tn��F�&e˸�֌�56�n��]SZ�
��f����n+�BRY�@!U�e��U��5K��PS�d�UYD2*f��Z�q��SX]l�kL�M����ShvƷi�Zn.å#SZ��+vc��8�E�i��i�.ҭ�Bʥ,xd6ɥ]�h֏p�M��A�4M��]a.����"j�6�&fJ�]���sn�Q�c�1�avn[FP�HN�H�(�����u��7s�m��.n�s�`F/N�r�ۼ���&�������v�g������>�U��x�ݛh�_i#��2��z���0Qd�i�lUƙ%���I<{�q�K�f���.�_v���km�9	T��:a&�e�e.�̗۽�"j��w
Z�l�@ ���x v S2t��������G@YUv �$�y�5��ݛ�uY�+"�������J���y<u����=��� {����F��A9������"�]}w����y�u��|>�ƫPI]���od*0U��C�zϠ�Y��1�:��ԤB&e^�:#��4kǅ�p[�>��Ֆ�Ki�V���e�ٽn�b8�^.�C"0��!b)�Fwh��fԠ>7T`"K�6�g���fKW0`m(6�!J$��7mE�����Y]��q]���m�i1���6�2D�AI�y�J�nTQlZ�a|�`TZ{�[u���<��a.�I�mRj���"��.�"��72��{[��wI�9���S��[H�(m3(8"1�+T$�+����z��Y��8k,�?/�����sR�C���psC��8�P�s��t���lj����b\7I0@4[%u�������(����җ�lY#5��T��4�t�k�pS8ܹ6��l�C;Kcd���֬�`ƒ��[�ͮi�ʊ��f)^���|���"�d��;���G��<#��&����b��5�F�j.��DMHq�{�1o�u:�e�ރ��ڤx32�8�MCO[��޳��O3��
P&����Ӻ�w���[��yz��]s��l&!���D�`�3b�:�#��Lʌ/�p}]
�0�DT��̄�7X��ym��f�X�=�y�}UΔVڇ �#�F��W
�v����ч�R���JU��DOr���z8�H�#g3k��Ⱥ�3q�"0��R�K���ۖɔ�����{�zȹ)���s+r�&(�oP������{Ù���h|FW.u���S�>��
�����,���N�w�qji�h�\���N�E�IM��;P��!�ob�5ˇ1�Ÿ��uI�T"�F}�@ ᤳ�z�ѩ��vD��]b�:�<��?^+��-��Dh)�M*$��lU���)i6��:�E�C SI���<��b� �Ϩ����M�"��A�P�]�f� �����WVr��j*��NH�W������3���(��T���Z�4ۑ2Q�L\�1C��0� ~� ���c�BF&E�����sk��� a@����Ӫ�A9$�Q����0&�;LD�u�=��p��Dqf��$D_]��7�oo`����Nɪβ�ig��ӛ�֭\*�gP�	�M&�1_�V
{<�<`�t� �m�E"I� �-!?8m6����\�c��TQ�q�����PB`��X�4ׂl�����=�cٵ�~���u@��5��"��s��x ���CE@�φs)U(�&T8;t���#΀H[�D�0!Yq/'����cK�����[wJ��>K2&�L����FƱ77���y.Oi(��`-�ro�Y�F��+���f�`�L��[�@Q!�JDb�+?��Sכ���܁7�y<��}���-)�8jx���?xy��_�=��!�`IZS5zp�=%�����^u���<Ñ2��R.`a필N�������h"�,����n�WX&��ٯ�:�?��������6%�OPn��2�����<�yP6��:����履���jǤIέ��}�6�+ao
�0�uٹB�6�2,�z+{o��-��2r;���j9�!S��C�����I�)�l�-T;�:�Ŋ^�;�ͤ����M����Y1	���o&NjN��Y�`xD���e�⏅lf�L�#C#2����{�K��>3�S�}����7��s/3m���M+0��p�Dy�x�F]0��Xq�JX�Ik��RO�f@{����rs�Y_j�3������30� (U �Dy6:ﷲ�bg��$�Gt�DD=bv,�q�S���o�~�UI��!do�A�������t�r��i��B��nli8����y�R�~�|H� ��3{�>$�J\908��NӎQ!�gՙ8����_6&qs�Z��1������=�@ qF����'ܖ>!����D����h@p����E�6bm��AN�����RX�+ٕ{����T���^�6k�b�J�9ͅ��fJ��2HU���U6ة��h�[U4sB�@&�v�mѶm�6�7��~�T�ݐaB˫�b��x ����IJ,��j�uٛ�0H�3 Ot�"Q�[w�N��wa
%	��/4�V�����I �{�j�������~�U,n�`&џdr'�a�tn$��M������Q��_D��6 1�f�V]����x� ��_}�*��)|��������?Nܝ�Wヮs�*��o!f�m���6��|���C�)d}R�2!�v�A��Q�l};lZ����q����}f����}d\���J��\���;ӮH�"�ydٞ�9�����^V�F��YI���2�B6}]�����}�^�M�tέ�h�є�mJa�-1���1��i-���>�����߻���u���^.ם�T�ef9�a���v�!Sl:'������5�YNl[�� �k��6v��g&����C�=���g�����`P��㫋��ř�>,�դNӓ*�tsݚNz�#H/<�H;Z\',��	;&������2N�S	ő.�B�@��.���S�P9��x�����g�{�U{Ц��עH��dY�@���q(i�7	�5Ԭu\�v���q$q|�cbμTQ�=��]Uv;b���F�hԤ ؇
A�r���j�q�*,J SQͻ�%Ŭb�z~���Y��vjl�r*y�BUP���(��tI�Sl����}�W��DwD(�.;;'4����^��#�T�ԙ{v�PEV��9��'�>#�� ����<��̪����i���-F=[�u@�ί{�ǀ���Er�3�K/#��{<�R�;pjk��-)�STi7S�չ�M�TZd|��gmv�Ԭ�#�>��\�~U���<Õ#p!���R�Ρ<cKz�}ؗa����ʦ5���\&[2��5wg�=�]w\�zn��JP�W.86S�=��ƚ}8y
�J�A��sB��P,���p������J���]��!���5w4m�d�i�uWR#��eUN����$]��CLS���Y9��]Bq���[�E6�qu]sz�GoJTI��b�ץ�#OtV�?d
����7Co��Xl6�iRujT��X����wXx�{��5�|��z��Y���h��Fh�!T�jZ�ZsSv�9�d���ۨ{�Nm�n�vf\�C^k)���n�L�d7TE[�?*��w�;r�����*�-"�Ff����Θ��2^���u�ޤ,���u��'p:�ղ�2�Km���%C���N�m�ȳ���}������E�CU/Vdi��L̥.��WF��֫q�$��Ym�6U��wB�Ħ�eL;$��ާ�2|y,�����*�!V qƐf�y[�u\ب��#� �wW������o�í3i�>�y~���7X�Wld��WS�/�y�~�����>�}&�r'�h��D�^Qf6�Y�6v���<6���[T���ƊQۚݔ�-�.��	�Y��F��n�cm�]���SWZ�*ɐ��{��z�oz�T���,��
��*
{��y�u����7�M�SZ�6欨�*0L8m�����l^ʣo������|����[:�,�+bi�Kd���фΫ�_M�v+G��O?�b�{OznV=ܫ����O\D�Rn`���c�)�����ȳ�ϥ��F�3ؾ_�XJM����Z.��:w$P��{�H�"&ؽ�Ż]~��	�5V���g��~U�����)Py�$����kt�i�EF&E�-��ܿ�sդ�z��Qj��d�j�ѻso���9=�u�]Jk��|�z�E� ���I���}�G�kZ�E�g�;�[;�_5oz�H��x,�#.$|�a�2D���1Rp	gKhV� ۰O�EW,�@���PvX�#h0�L�~YZ4*�V����[l���mWl����
�vV�V�"خuX@�����̯8UW;�i�R��� �{d>  ��� �@ ��=��2�X��xPk�Ъ��ww`�$t��݄�����  n�����X�PU����/�E�-����nΛD���L���Չ�C&�ݡ���1��.h:7@W%���J6��4�.Bۇ*sJk�VgP����-�cnRٕ�U�����*�F���� �KP��m5l���c����ka�,0,��ƕeK�������fղ��B�L�Z1�%f��"�]e�3aƶ��*���e!��J������^��|��z͊U'j��2��O�L"�)0�7%3*sH���(�|��T�B��Ӡnm�v�3�����Gww[�üKI��۠M�C}�ۄ��z���.XGnV|�fNӀǬ�LL�k��ʑ�g5K-'k�A(��"� +��0B��0�6K��x/Hݒgs2"5��m*�vd��p� � ��{�x aҩ���� J�z��T**����{�������Q(��M��j׹{&d�q"l=�_Pm�g;!��!��K
�����43��YMNc������7��v5��[�Րt8l�������D��l-��wa.�{����G��o����$q��B��[8 |T4���{V�E(�E�}k�rs����k:�7��j���(|�n{�g|~�$�eәq�h�!nk�$az��O���U�@�}����q�#m�����+����3��{<��"�����<��J��p d�.	Q�EA�vb#}X�8H����.̎�$1��T�E�[]����[WƐ����Z��Cj53�T���K*	�H �S!��7�ݬ��WǴ��Gcb�,����O3s�7�&.u#7�	s�����W[�������4i�B��OV0�$1Ic���d&BD fYI�Z��\U� ҍ(Y0:& �I�$���;�1�%�w]��0�7�d虈��{��)�fw���@�/xx.j=�hI*%�ڎ%��>� �b{7� ��0��jVCZ4zj���oR����z��m�[u�Ud���0F9Ku5�|{z������2�!Z -S]F�
5��kCf�*�)�#Oy���&���Hip[n��d���Ïpi(�i|�������a/Q��3;�{�5酤X��j�y$2g1��z�laW�a9�B�=����n��J.��`u�����<��W6>����Oȳ��7z߬��1���/��љ\E+���p�Dy�N]|�_=����>D�"4(�8���.@�7������C}�_M��9wyj�3��S�������@����6ԛ�^�ʈ��C�%�T8�7.��W�[���eK��AV(�R��Y���_g]wuVMbFaB::}1�W�>��u4��1h��^I�G�EەA�h���Il���֪��+e������=W��ĕ�<���%D3���l���ٹ�\|5��ϕ�6c
x��>=�N�vnU�#!�5�=��K�,�wg��S�٘Fm	"l��0�Bͪ����j����"�ӕ�� �<�;��Q��o���B����@�̡<�w�v)�s��z:j�ۆG=D�60��b`B�Di��2l��Gb����y~��^��6�D��}�����8�ƘLc���[+qb�v�ggZ��0\�1�5p�56�<�L
4�٬�dw5ۛ��V�:��=�Ϻ��ŗMҘ��F��D�� h[w�~7J���@�0�lSFJ�����[�����z�YzՔb0���A߽���?�E��]q�=\���Qk#](k�x����Y@:, �%*o�?��̣�o�AY�Q�����E�.ss���׵�^�k�Z�#�WbJ7TEX�=��omVm��< �Z�o�q~�c�x�&��T�������Φ�����LY���;����DV�cٻZI��$̖-@4궻#rы:�$���!es����W�T�W.!5�QN�:9���	�o[��u�\��\���nQL!��uk)Gd!Y�/%b����(��u7�w�'���&,'	2�)")��6�������-x�RH��m��9U"�H4�-���ڸ�SJ��i�)������r�1�N�*7kBZi�N��{�/]8�҄%9���N�-����|g�6S'`I��l��mA�Β���i���rxb�"��9��ΛvD�:ӡ��DU`�>:���ޛEͭT�A�̲d]����D_G��H���DB�&��=֫l36�0�ʠQ��轄d�d��7Deb�{h}�<>Uw��ϭh�㪶q$7J5]v�]U��;��5vu����R	���vmĴ��*�����v0�̊"oU�t�Fo.2R�����4m�E���z��w�&ϧ;��1�
-���%��M�f��x�-}��$0��jVCZ7�Y���Ym�����fy�!���/R�Y�l�@��{Ç��f�pf���$D�a���kEtM�u��7[���ae�ܰ!��~�$�6ƐegU��gJ�,_[����8�Ҕ�ZW��f��v�/j'`#Gd@��̞�I� 's�B�����)�~�:�*�&ЀV���]�y��MVڿ�~�o��'���y� ]�0r��T&�L������R$�!~$�Lv���n,�Ϲy쮨������}}��+/b�����0
�7�Lyј�S3'n�z��ެ��\}��AY����w�v��l�WSY,D��ٸ����o�Tb���4䪪xT�D�(�8�8��L<I �`@�[
{�snwq3O+1�\M�E켈�7f%�<��xxG� �}��'v4��W��HY�"7�˥�&B�rΟ�
��������8�d������d_�eR�{w,�T�%.$[���dM��o� ����B
	���I����1ȍ>=��0��7��!w��Cz�ⵊ2��
d�f����[��AD�
���\^N�tk�qA���NR�j��@
>��ݗ�n�tI��$n�$VA�����J؍&ܠ�����)���23�".r��7WL�ٚ�D��ۮaDئ�����rw�!��װ�N�d��V�޵� G��S�B-��E"K�sI�Ym�|�������� �g�����Զ��k5���*ܰn͗�صh[uRƪ�i)��K+V��4� :[�-�l��q�%؀,6T� HA��������U�9��VdLo�����o�u� �bX��M��[�~'w���߈��W:㖍B@�4�k���}��wg��u}�ß��������!:�N���/K��d�oU��O H��҅8��a��;�x{�s}�hm��:m"�T0�dq6Ҷ�F���Bߟ�+Kf�ǀ�Imԓ]27�xӈ���,b��^�"tƜ�PC�ެ��Y���A�LM�Kej�	�!2:.�����im���A�kH�'N!X ^d�0��Ѭu#��Rѩ@U�y��䪍�5�0��6�2b<�]�Q=����z��=F�PE���P}6/�:dqe�)){�Xd���6����?~���]w�^.��5����]A��jV���K�Ŧ�Qw��Hv��j 4�"�ޓw��9���v[v��V@�8eӚ�LD��1��u��\d���5��dc1�1�fvq��: i�sF-��)H��ɑ�ק�T��ݱG�:�Y>dm�ֽg�P��巽�B��/RFͱ��d�EV ���f�����Zo�ytu@�Z�I�.T�m��R)V���
�G���tA�6*a�3�����ʴV��ܧ��h��N���N�\7"��B�$�iC�����e��h��E��/e����᳂�7�y�d�Q*���`2M�If�\5�i��N��!P}�������[c<�t���Yf7,8���z�+��	/����30ey%���<�jK3��.odx��Y�������cSÕ^ѯN���ǭ\V�ɵ�8
B"�����"�&N�c��ʎ$*�>|��nurE�+�T&�v�|>��������D}�$��N�1��.����f>��l&�s�?�������޼�06pk�r���A(a�4���>dv@��~�y�])��{���P���-�l���ޝ��j��1�d��2c�"�WCw�9ϗ�fY����̖-*��wuDU�Α!'�,��lfƙ/#���[Ԅ(�����'�V�NEIҵ����S��w��@h~HnU��3�T%�I��3Di4�)k2��3(�؆�Sr)�1-�����E���l�,��F�J���C�RD��0��2���	BX:���f5����1�x����IЬ�
,�bo:�!��7l"�s�� ���(�
!5�`lH {��:������;�����m�vͼQ6�H��!��9�v�͹�s�Fօ��@CGm�]�s��U�W5
cG9�s�6�U�v�-L�s��m��m����;l�9�dLͶs�\溰��	��*.=�f�s32�ot������=� ~������� �H$��32���I&�� ���N}���$K�R� t��@��  �����;�9�<> �S�v���stL%�lh��ٵ�.��	t��kiW@���j�k�N 0Z3Q)�j�ԍ�j��.*�p�c b�B��I]f�l�x�0q!��v1�(�Yv�C�̮ի6�l�nZl�i����.��&�Zf��"��؃���+1[Q"�l��vt���̦4�Iv�&��CP�P����-��W�<�%1n��ۭ��ԻF��ئ�MIm&"9
���cgiMq[[l%�!��� �mZ�[Ja����Ѱ�/0��(��c ̶-�6B:eѥ�U	K�0��Yk��i���J�X��h ��$*�3P�m9"��,c��%д[�8��t3�a�K����җ��鳛��ݻI��P��ww.��#yw6�{ze-{�`����v,���%�dK���Vl��˅3%��4��fU�9��A#9+ Ӎ2JX@eލd�ю$;D��}rQ�����TY-]�p���VA�h$s/.qm����u��mYz�`�d���I G��=����G�oB�胐@֔C�)�x �g`wzu�������T�m��	�=��X��q�����}U�xD�̏xx}=�(��ڏ��{|+��J��F���(٘ji>-�DI�E�ñ��2��A�Û�!Q)�q����}nU�mS�l��|�.�!M�yMX����ߙN��'S|��F�-J������U,���
¨	�ሏ$߯����8��ݍ0x�ؘ`���9Dm��i�nxy�ە�sJ�X�$�ݬ}��o�w:~�#\�C]�L�����]��L�T��4d��_G�������)D�,QӾ>���U��KP�m�d���;�� ��0��[\w`Iz����{ʍظ�m1h9JL)�-bl���0�D�޻���%%�"��9[q@�����&J%RP����b�o:�8��\:�i16��%[V��[�hZ� Sk��fh߾���/�<���[j)ζg�{����Wy�1����~�5�R3`]Po�|`��w݄;wLۥ�f:��ZѢo�o�5O��%�q��#���;�5��#f�����)6��c��5�u��۬N�Yi�[O9|�2�:w̋���?f��\�0dFU�\����w�p�ʂ$��G,�Z���y�b\�T�bHL���,��z��>�O������ܨ�U.�xaj��;���dl�jZ5(
�^h��ˇ�/Ɂ�.8�_j�U^r'ΆZ'�-�1s$"�1}�?��� w;��S���Xh%���"n"�v�DX��;�� iߣ|���tk���؂_`��弒�����vp�5������<����#��}���դ	�����\�)�i���P����hT,�VC�:�}�ߞ���޻�3ߍ��	�rsߗx� ˴�\nl�ʊ�g�Z^��b��q��d��רo|=���/����рFU��
*�5.�dnZ!o�O�̻X���i���v/��Y*L�{M���{(0�>*9TJ��فDE�b�7�r�2�zwdt�+}��!���#������\�:��#�OF��>������gV�z���q���Wf�->:���(^!X=:�Z��im�h1�w�����EI�kAEG&oe����&
� �CSQ��9�q��1g:y� H�A�'N/���'/$��P�g*5t��4�4�H�(�o��>�H{�x���r�!r��ٕ[y�9��Y���sVҷ����x{۱sY�{�l��+>F�M��	)�u��	M4%Xv��ADR��[��mx�G���^�ӬA�ܔ��y�!4bfD��ݡUW=���cNti�������;�y�<���j���^���_��%�$���EV:��-��N��]t-��m��3Y�j��}�*�"�T��^Ή�Q�g��7�n��=`��f2w�]O�������L
"2��fK�_{���w{���'��P�>��F��5(&/�����ݓ^i��]F��/��+�s;y�*�b)P�
7*٭��:x�׃5��gh�m��4�-����U�
�ɷ�1ow�� ������o���kEn$�kT�����Q1T�;��=�LqA��思:�h��Mu^�4k���v!sI�%AD��\Y� K�y�Uk�-�:k�ݶ3Eq9�;�NB"���*#�$|�_jr���Qf^9R�����E�O�]�9�$:Ϙߡ��y��-޽��DI�tPU� �s
I!����_7�u~�.^�q��p|�㻫�=f�ګ�{Y����Z��f�	��wj=B��r����ۦڃ����k,��|8ԑ�lI�.���ND�\��#m�=d���[�N�?�������s}v��� ݌���HYX@��c]G����^v��t�}>{�����[in��45��5���vQ�Ů���ڱ��ivT��36�����n��y���+����ex�E�nwwҸ���UDD��� �z����ʛ��8��Pƹ��j(�f�3G�7κ���-STC@���8��N��I6�3��ʐ��'\�>�9b��?n��\�08a���������7�/|3�a]t���B��i����?n����;�A}#�"����(1D�i��c&g+��m���/ �8Z� m��Df�<�*T�HYk�p�X�'�x�_E�5@Ϣ��'�����#�PeH�f('SU��|:f�ۄF3��la��~&���q���RF-��-�C�9]�}�g����feX5�lz�-�t�93�0���ݡ��6~�Zx��^�z`�q�
��~�@����0²��l��1�k9|�[o{m<J��V�����]D�~{:�K|��6����.SGWkEf�Q-��)� ��X�Z(�� �%��ݫ��uʸ{��u��0���z�{���MbZ��U���Y����>����"�W9���]B�TGTj�	�Y-K����Գ��ooB*�7[g��Ʀ�v�O*�M���7>��]wI�V�����]!D[�V�swrwI[�O���Rv#ۗ�92`����vk���w�ɽ��wGWE�p���F�/9s3���U�jG���-ʰ,��O:�wJ�!�2G�T6f�d@x[��������IחүH�N8��'Z�i[a��D�~-%�"f`P�,�������ؒj��bF�\Gl�}�z44ёƦ(wD�����9���D.I+ۻ����Cvv47z���M$�3���<<G�{����v��dp�^c#l��vr�lW�u�M��q�
BɈ�����i�}i�8#'3e��T�����B��{�uG�bMF�k��]�<��A�+#7PDVb��z&�sw\��/c�/��wUb��:�5b�%KE|��B����E�i�V�o���;d��"oV�=�,��p�r��K��*$[i���"@����.�Q
-2+c	�ͼ���q���������B�(ܫf�M�u�������q�����7�x ��ŋ�����e�Bh�y�1�	�l"��h\��� ��(����nkF�m�ov��j�.�*j�NÓ�3��kos� �����  ]�ܩ�[��|��Ӵ���l��X�)*�޼j���+Rd�")�+�벭!��4[r�.��r�����B��%���˖)�S�����1��ҹ��}�����dIdo��{�w]z�{���m�	}�}�c*�^o9�7�ƻ���#�n���/�yW��-C�؊9EF��Wj���5��q5�2.�Rs�j�����ij���W#�R؂ꈥyμ�Q�؝����2Ntiqًz��;b9ע�]ڴ�W+E�Ǜ�S�خ$����/1������[#b�;a�K�g�=�;>��~+��={��~�v2�9�].���D҅!����(0�����HMY��i�k�`Yui�d��R��3v�k	�%�neh����=$ѻv��˻�~���� ����\��s"��f��8�2�R�����#O��FQh�H 	�va@%O�~����=���O}�{g���}�z���=t�:��Pl��I�4I[�LaA��*�i[:Ր<84X��u�n�L�.4$(�9��kr�3�3I��$-Ԉ��
� .�7�IU���J��Q����/���R"�/����~��;ێK#`Ԍ��Ar��(e����d'x�D��O�w#zׯT��_n�z`&�6�7iѵE�2�ʬA���h�a�Yk��k�u+n
�'�|�����Rob�]P0�/`���M�Ď@2B��A�&����كEM�|I�� |-�7ed�h��]S�8,�27'0lH�P�{�j��Wz�:��CoF�e6@hy�6(m8���0"F����>��8N&Eba%-�L:�ѷ#����ca	C�u5�XL1���>k�Kg:��ԛYy�w~?� rЪ�6��u�b6��v�mT(�� V���V�I�,U�m�\�Q�k\(��l�f� )�7w` �H =�&�u������xP���6����$�X��.����� �݀�� �@����|�3��W3DR�5ʶ��)ɶ��b��3E�-���mwP�im�tu��,5�ݨ����k��)��i��U�*�mf�Uu�f��הd��pYF�-�jM-h�ڊ�c���u�,��s)[�-�P�gJ�h�ض9],U���7�p��Fɦm6ήdl�qR�JQi�u�U�іe`ff9+�wS͎���4�w.�e�9<��ydo��L
��@�u����ן}ߡ��&!��
a�"q�n���n�3z1���o�t�8��q lNU��<�(� .wZ����-oV�� ��VkW]����$���+�Ō�)�)$�>-&���=��d���ڻggv��kn]�wF�+���pQ�{G����g������N:��9$���rFw{���b�,+Ch�t�Y�S�j�ܥ�t����C
$Ch�S3��BV�+B[3��A��rl��f�%:����o{�}i�9��^�ݜ�Z�fϰE�P8���-�e�$��N�{cr�������־�}����F���ko�p���B����}3#L�Aj��"Og!��y��.120��OI؄�[^����&L̕�k����Y��6��vw�r���DTrf�PɞH�BZP�, {��.�xUJ�̊�Õf�3vz�1U����YmQ�کDU�~�^�#²��j��(�E�R����)���3�OD���"�Q�z����ЛJG?��1/�؇(�$4I(�O~���ğނ���d`/�0v����k6Fq��ܔF���	0��)��^������ {�<|��0�"w�-f^
~��eխ�xӾg�w���C��T��U`Q{�jf��ν�̍�Cz׬�jZ���������K�L��Ń�P�'�t��bM)���E���!��I!B��wT�8�=�n�|{�ӂؽ7�~�� �ߧs�{�Bȭ�
)2���d��*ˣb���V2K��`ġ��Ka؆���㯬���[ׇ�G/6�wt�*e�f��$m����Q^�n�޽�~������^��8��k����I�ւ0jS2��-J�%F�{�noO[�4T�. 	�Y�uT���e;��t�[�h�H�"O�H��2v>�a��������M���Y1���E����U����������;a�j*!o(>ɱ��!���'QV����켼�z����">}�lan����Pw���DV��&S�*��^o��7��hQ�ቭ�l�Ĩ��x2�W��G̎8o6߬��FǉFt��e(��S��OK���x!j��Y�Q��g{�.�t7\k�a5QQ +;�L��Q�bh��G���������gѤ7��չ? Ss��!Dl0��d̪)*�"M�t"���#� <omv}�Jt��Hˆw佹x�F�L�F�{������G�>+�>���[g�/뭽m�:0j���Ԕ#G77M06���~��m�Zs�}��B�~2��gSWm:-t%涕�BR�&�1WKp6gZ˯��-�p�ño�]�T�u�04ns���HUy�|�����݈��o&�E
n����3����G�����3)Y����ȧ2�!L�4J�;��a����7`�D$N��	�j&�
AטP�����?����u;ʯ�Ҧ/�V��9.�.��q�J6�W�ӗ��G]{� ֦NĐ�Ӻ����`��G`ĊWh�Ewkn'r��ݔ�b�K���>��;%����b1�䌖�Ar�w+ד�Q΍2��"%>�F.4�b���U��z�6Qn�05�r������I�_cӄI���ş�n~�~ۘN���'�4Z�e�Ԣ*�φ��z�Ժ:�3�[��Zl�,1*����<.���~���"��ɘ127��N��;�G5ɵe�_~뷪��ܼ��U���pЩ�J0�,�[q��6���S\�.�B�l�����k��r�v^kZ�7�gu�WH�@����o�~�kv����QE�z�ί��'����dN��_.̬͝�"�e�����(rd�jJ�5�ߗ��뾣�$+�>�˹�,��L�� �)߷s)EJ3
S�Q���1�	_w���)�Ux@�1�bx��\�⨐���+��VfY�q�����Ũ�MUj�� >��Z�eJ𻸆�R���O}���(�i�a�����8]�q�cL���}�{%"-^�@1:�� �$%3��X�����xn��ۏWm1&�8��d��^k	Ӻ�=ڴ�@3vV�/ʌD)��ً��=�?IO��Êb��t��bhaf��� ��$�I�� ��Kt	� �0N�������@��٢f9�a`:Z�"�E@�1��<	�>��LD>����U��[a刕�c�{�TM[߇� #��@�}3'�s{��Ȭ�7l���N��{b�3��a��QU�:⏣-�8~�����e�z��~B��i��+��JӢ@�V}�z۵�(X�N�Uф���2�spq��p}ݱ�Y� �K�Xb�G�¶����e@&�|�"\thk�Y�[R����_߹��[y{�֊�$��4�㮝�He%bB@� \�c�z�,O���>�4�"���N�^S��%�6�>��:[-�t�$"(�=��r������:R`�D*�F�M��Q)һ=��lʲS�z��-����j<�g#�4 RD�D�$�&H�%�g������v7M��v�b.�ӻ��\�-�{������޻�z̼��}׈nJDV��&S�*ᛁ��𺼿���lqϣMl�Dx���~���ݖ��q ��r�	jJLJ�r�~��z}��(զ��.�!P���{�=��PU�)��{���Y?,�Ƥq�I��I��0�om=6M�o&�X�}���d7�����y�����ȹ�,��P௦�&eQIT�oyY�}� ����
5���x>��a|H�y���bd�Q.KV����e�ь����u��qVm�Z1;z�,���	� NJ�TS]��1�	w6����Lx �{����b�r����D�M� �knR픓��Da9{po�)��j�In��b��������b�r��l.٪Z��ڭ,���T���m�&��rj͆W^m4JJ�>{�}Ocv�v�mE9�({�����w���κ�9.�B�V*����
���S ��V
в�Z/(�2\�wr�Y� �ب����|,i�~�7]���XsF-�o�-��{���^Fv.(�}�law�Z�}'�v˒1nH�pa��7�����{���\q�������g�o��*����Ƃ"�m�QP�Աb�X-��$�����4��]0��/r��Y5�:�4Z�,��V_{ҽ&����]������˽�o��ξ�^y����2WY�f╀3}�DT����2��"�0�A�	L8��K)goL	�,��j=$m�����=���Zn�W��W	�A?a�{��3%��a���:(4�4r���YSbR�.�R��)�y��e+�0�6�������=�0���w��A��_yix��Xm�M�����Ϩ�6�qB4�D�}��_��}۵�H�|���Q�R0$K�:���ok���AEZ���K��G��]j��TlZBV)�y���0��뺊Ѫ�TE��=s�9�	dZ��������}�����k:��ř{���Vt���JJ#oAI���"��xjq�x�K�P4��۴ڒ�z� U��{�������ޞ6}g�vDD啚K��>�r�=d ѕA���wh�l=Bq�j�;cv�DVFq��݌�d+�G�5��5
R3S$�[�C��  I�C L0�iF!�\�^y�}ff�kZ�ˬ��Q�s��ђw2�\�s�� ��R{�M�4x��TD�v�}vro�r�1�V)X�]�$V����t(��������9�zH��B={���U�b��ys7��0�q�����yV'����=.�eԈ�E1F�5�����	��h��T�0a�/�hbZ��\����;�����'^m�������g�t�̃�|����n1��7�jf"�D����x��LF�B�X��H�Vc�%G�ot�-Ď�U(�����g<9W۹�G��9�/V����鏽�{�;7��2��8�.8@�0����7�y*�Q��
'�� ��є���qu�3�!�K�H�K���OR�o|��x��bQ�9fM���ʌ ��:s��B��adE�����������2"ppĲ�^I<���7����o�l1Eαg9�s��t@3�&���4��q��ݰ!��s�.s���F��Wg9��ttv���u��qC!�ֹ�m�����u���9�v�; 9�]�s�3sBۉ�m�y������r;��Cwvܒ �@ �Hs�%ə��zI$��� fHg$��K�I�]ɹU�.I\�I`�$���*�NrL�ҪԺ� ���R���6�Cl�Uܘ�j,3J�Q��V�7ۮnf��*����h�M��V$��6%-���6٦��Y�:�ša���ך;V�%�K���*�?^�N����t�%e�+�-�����%�Wi�L�0�q���@�1ڎ��e���������	.],j�]��ۊ�60ۜ�]Cg5.�WlK,���(�g-�!tunXLf���1�l�\�Cm].�5�kZ:�Ѯ�3W�Cm��k\X�.Fk�m�Sn�6:�c],�E9�s4�b(-��ٵ�h��ସ�\���U�siZ��̵
����9�� ��ZL�6�6�O��T,�YQ۬n�ش�m���n���V�04^���-nTj���]������-�A�%$S)K��ρ��U��	9�B���l�7r�gs����]$�@�r8Im"�{y��K3��,ly�6q���5{w��a�ܱ0!����s�v���ՙ�{��I6��n���J�� <����������m�B��(��K� 11��M��=Q �	�К�T�|�u���׾��!��/���nK�P_5��};*�w[�P�~����9�]w�{�O�`��v:�Y�J��ј���̍3����z�I}Y���#/�i��5[���K�8�����݁r��R�K�z�En쎄��4�R�av.ɸ�̕�H�����Zg�Ⱦ�
�\"�P��(��*TK�=�{�wBK�`3�Q@��8r������oo��yڴ~��@� ̑(ԸE`�u����� �c1�I�Fk0�1n�Tָ����S����*�����ªP;�ئ���*p>����7+]z����b))�޼f�QF��I���(�g)劣�LC˱�\Se�Z���L�C���Z}����.��g*-.�&��ukq�e�5J�0��ӖTH�؀��fЖ^lc�E)Eó��m/:��YaSY�Q��b�?���}���0 M�n���!��T�~J*#�;FW��m+7Q�ر���b�b��aP�k���޴�;f��a��Q�i����`��|��}ǫ9ɒ1��.����":,��h��v�6��?��8���ܪ#��gr��؟i�������*�P�?k��Z����ή>�昣�H��N?���:�z����.TZ'�� ����ʬ|�����;3v���[��l`������2W �����St��b��8�~-z��)m�G����`&e݊�o�{��_��:'�abztuM�Q���&j��-þ��1ȍ>���聄�r��o��5^�3���b)8I��]�|��C
��ty��s���}/~k~]�(hA�Ur�m���U���CA�Э���L�H(ewu���7e���gwF�*��e��u�M�f�,]�U	�*(\)Ɯ�Tx�"#�Pg�F7�ت$�,1�=���eF��`b�o?
��ݽ��	�aa��D^ED+��/:��tbW�V܁�>^��| �`�G/��TA6A���VwT$�L�b1t�5׹;�7Bfǰ菗�}O�ޞ6}z�n����ZE��װW�R���z�K���ί?%ۮ��;G�!tQ���
!�i�ӧL�w�j4���uo�P��&���@Q�2w��"o_M�Z�*K*8�q=� �]�ݡ���:b͑�Ӆ�F����k�3.���k�	!dI#�<������e�D.��}wv�3<� �;��/V�S���� LMkd\j�ƒ�̏Iq����}u����X����d�"�7��m�ᕦ
y�����f�\��t��_
�lE�2�&*��{��U�w�ۥ'���X�O���Z ����1U����z�t�܆����}��
R�Į���TA��H��2IKe�����P<Yu"/���b,V�� Kr�"j�Fx�&�i�m��w\�^G��[�ő����Ś�Y����m<AuO�	_A���D�R�T����?{�������ϕ�x=��q�;�����k�ߴ}�R*b!�N}s�TD�q��L��ki-�X�m�owTպ�˜�7u{+"-�ى�[�#� yQ®;�q�4����b�z9E]�,[�+�U}_TR]����h��WK����տ{�Voӹӽ�a�/|t.��w)����t,T����&�:y��V�㵻:�F����:�Q��'�NG��+�k�^^"Lhj\�:����I���s{��߻���#�D�lf�?g:�ϖ�#�o���^0��'"E(ӯW��  �~��ǀp-Z���w�Nx��.��%�O��4ʇ�B��E�\Y�2�1r���RR͓�y+k9�ҽ�f��"��5��#��,�|�tan֐�{�IJ!
Q�
����ݬ5�o &�C7��-Z���Y�^��H�%}�3��l��(��`����*��si�
hMM�.v�&hk�\�!�*:�[a�j9��� ����I�5�B�Q]��R��~����v�w�J�בJe1c�x�]<����ZQCF@�m��p�]E���P�}eU������q�1a�m��ĮbUO�{��/5mǬ�Gh�"-�hp��-�&�IR��'S���^���3�&J�$����Yw:�=h�#�4��U��"�pBqK
��i~K~���k��Ho1�sV�wE�s����1&L��J[�1�{MбZҦ3���zm��?AZ�μ��ٴ��@N+�w���R�2�q��'��#�xr������c���+�.&�4]Z:;�V=d�wXӽ}C���
cWb��4��&se�OU�}4cn4��ZL�ر�w������6av:��:�n8�{��u��1-�����]$�2�%�q�5sn�
Kf��h#�1�� p� �֥<�ÿ~ǿ|h}�뫚;�'e*�/�H"b�X/`�!5��Yc��,�����N��ˮ@�P��A�����.��2�g�s���/{p�م�.4��D����y����A&d$�\yo`��Iލ3Ҹ�>�TF�.���;���kO�`��C%����MxT{��H��܌�Zlӧݝ�)3��j�&��&Ud��F�\,}���m�ˡv�n\��R�C?~�����7���d���.��|+���^R�\�X��(4\�KJygw������Fkc	Mw���}}����d^�:$�wuq3���Da���� ���]�I;֗�"˼������3��|��9����^N���lLI}g7��,�ţ�uڂ`b$_�gGO- H;������n�ݢ��N�6TZdWс��)�%�$*}��Uf`�z�x���|Yb�������B���"��^:&^�>#w�� �b_"�Bе�]�YJ�Z���}�<�������� ��Z�H��64D�%���b��%#�6�t�ْcGz��ܪ��E���3dw fn����������@�1�M��i�l\�uLN�u���=6p�Z��y�xp���eJ3��te�&�q-4|�k��x��G�T0���p��Z�����Z�ݖ�LB�6��_]i]���:�z�?P�w�Wn_�-n@}�Y�0�!�6%�m�hh�=�)z����c<t�k�����k�;G������<~E�2�b�
�|g�u���ʀ"h �0�,R�AjM���x�g{��~�N�:�z�<��'�C6��7��tՔA$�B��.����r�8^���XƔ}'5d�`�$�Q���L�0�Ԡj}DVGw!ʧ�7ot��a�DQv`f�9�TR}wվ`/J�nl�-r���~�}������oL�� ���cJ#*�t��j�R�Z�W//����7ǅ�~u�M��^�����4R%,����nn�=�hʪ���1�b���ߞ�����5��ߟz�a	�� �勉�Gqt!iFWwi�������X�Ͱ��l�mn�.!i�al7,.��Lf��}��{~����BQUS��z�/z�m�g�[���}�Īd�#ōq`���$��fH��3;���nӢ�3bX�_߿~߿�}��s��]ʍ�k�QH���i�P��@:d���w4�V�{X�G�c.^�!��Ү�7q���,��}$ə���/Hdfv3�{���,p� y�A^�����t�FQ����+D~��֜����������Y�Q܏D��)s�6BE�aUɮ��ϖ�$d#��MF�����zy��T��k1�.©�F)@�Qcw���]=C���Xs#�s^b�x������d-Ԉۈ���qc�hR:��	F�P`G ����>	E�bŴ�ɳÐ�e�G��G6�\�bB ���;�7&��%�!�R��:�Bǥ�nr�f궽� �Y��i�� #{��B$`%e$V�!�m&8�j���#$���b�ŭedMڏ�H�
y��vpr�{6�
��}�,�U�\��Y�H�)d�o�e������F�*��UZ�x`ͫ��r]fVܮ�\j[�2�PUmU�inF�ĕ�W�s��̀��>  �݀I  �$���W{��� � w�VfzK�]ܓ�n��O{�~��I?��� w�m�݀UPw��ߕ��I�d�.8��Ű�H�KF�M�c��F�m�YL�N7R]x�aJ]Nb�F��edS���[+��t&�l�e�%�ׁ�Km��nm��N�z[n��X��SWQ�Mpk�Y���f�6��v��7��/ḰФe��:V���S��*�	i��ͤ����&��6x�WK��s3k,Y���h��h��M��Yy
�e�!=/5��j������L�B�Qz��כ��F������d� �m`n�w�{u4r�����ۼ��$=�z$��:o870w#�z�l:��[�V,軼�Ni��n���,�Ih�-�\t��PC,���Ӄ�5�V��uniZ��椓m�JU�*3tE����{����BU ����⦀5�XTXO�#(qQq�WJ� 0S�����Z�٘�L��D� b��j��s0�m��7��e="�3f�`����sk�;Y��c`#tҶ�5H���7xЈ��G^JE��x!� Wӳw�����ǽ�����o��''x@����@���5���f���AB���(V��fT"��xk	�=��k��Y��r��g�E��tkj�/7q�f�
�Jp��j�3ӨI�v�t�fmךssf�]ʎkViQH�rð+/��[(�,��]o�E^����]���n��5�#TT��X(YE��h��n,q��"b?P�Lx�/�AMC�n7{��?l�q�H��vD#sZ:�)r��d�'&��������/���9��m��=�����k��ގ�dĖY���b�����זI\���n�6���z͒Y��v�/E�p�ܫ�����Q;I��W�0G����S;Ն4oO��j2T��Q��}im���]�P��#^�6k:Pa� �yW�,
M:���*f�E�������A�������(3,�m� �����q��xj܄�=�,����8�D�T'��DA)4a1ٽ�-���3z��Y�a�{�A���Y�Ns�X���b���J����d��}�scY��S{�z�>W�/����Y�vʎȩt{c�34��of�)�17ۓ���ᵗ��d�(��.X*��?~�wVQ<����M�a9��I3DA��2`�f���t�nk�s��f�f훻��U�Ud���׳~���uV���=��p����9qCv��^>�u]�,��
�����7��|�gY�@�؅H�]�碤�������2�J���P�ls}]T���&�2�#������@��{����!��a��J�����z�?#����ɣ�VwJ-O#vA�k���ɗ���k}`�:�S��8	��W73{�M�H��R2�Z�ߗC�����w�?Z�k�e;o�T@�n���z�g7�
���P�铰�����Ճ�2�% �l�T-0;:`��nv?u�y�O�� ��O�>�r��~4�̥a�L,6f��ĵ�/+XTl�+-�̬�-iD���+mfR����봤.�BZ����%�Qt(�h�q7q%�Bkl<<,9̝��s�pw`d��(���U�o�U�/���6�F�tCh���&">I&�e���o�ܝ�V|��k��^���a:����M[����[x�����t*0��e��yB����.+[�t�G�
P�w�z�og����|����쇖c��33���Ӎ��:\�z�#!n�~5�^d���8�&or���r�R�+�w�|��h�Ο3���K����|�)�Wqڦ�1G��f�]�
;���m�H%>a��-�v��pu�Ӯ����������t��WQ�0��n$��RSP�%boqI�M*�6�r�V�֖�L�U���1��R�k���ѕ�u�^Ͼ;�W:Y�9VpP�j7UU�0����6��t��|.Ǟ|q��{ܣ�ϵv�|<�s�������g�J-D&E�	��[��C�f�i�}�s�������/NTB���-�"����b������gl�^=�{o�Mx�F��:�;�3ޏ��昛�/K�~ {Χ��2:��V�u��T�"f*���zFP���To��-l�&@�
��T��$�����q'���z*�mu�{�?O���n��z�k2��j�Fj�k�xD���D��oeT��S������X�����}P�]�J�K{2���Z&H�D���4{�l��3��{ʪ�s���Lk�0ҷ�T�o��n/�nySVU���g����������|��6L�gȚ�ҐQ�%ˉQ3q�y;��^:��V�����������p=7�����L:6��?$������#5B�%�)��Js0��2���;܈��s��?�P�?=��)��D��B�Yd�w��d�ąB3�QX�w"�sk/�}�����B��p���=��t������oq�]��pD�v���B��m�9�oz<�{�Խ�JE
�,Oyߟ��]�m��t��ov�]�b�\��[٪�� {<�f��5��1Y(t�s���m� i�T����V;��Y��P�÷!�=�r�gWF��,�qU�V/O�����t�g�RKt�Y&�/@a�A��W|����s���4��S}�~�����w�l�:<']u�K���̋[̈�ڝQ�bKj^��������<��y_�G���3���u��_Z罬wZ�{�eu;�͊}�%(%#!�n���Y���ꉼ��/y^zkH�D�kV,ݏ�}�W�Iv2��J�S���3�[wd
���5�7c�D������(W�w���x�%�]�oT~DҢYm��Rm�#�M�)̲�,5�B�xܮ�\L��4��3)�[a�i�[��P��LRa���}�e�&��n�K��TM��8 �}�ӝ�l^�e�<�mT��w��Y�2�T�d\5%�Z��Y�\���o�{|��uソ�S����)��O�_�H�VH�a�I4ۆ�ܜ|��V�)"���+yK���;>G�jE.m��h�\�g��t�;-!t����0{\'w�����e�@�2�.���|��c���̡v-/pPa��=Jz�0լ9L{/&�wV��ґc�;�pN�JMr�]��F�f	@'6���{�R�$�\�m��V�<F�A����n�سf��::���.�W��La� ��R)x&�޹׊�dK`�������^9����MkV�a�K�se��b�  C%�j�ssp��3�\���O%T�� �x���+������y�-n����޾�Y�uV�k�;o6Fn��U�ma{����w��5�;�ȥu�]̵�V�'�*�����Vۙ����pjbqEvA)�,�����ٛ��;����[羔���C�F5D�n����˱�\�f�\yl��;��j�^8���l�-!wz�޷���!�T@O�(�T"b
^����Pa���-u��s��bvS��,�I�9x��j�Bm~I��󼿽\%�# ���:μ���iKФ�_GZsͨjm]�T��
����&<D�-ff|���˰�+U{/#6B�V��~����r��C,V*ަuO/qrw<���#tc��L/����V���O�Twl��gsp:;�8�аc��=��ookq?8+��po��an�����Ƴ�.˜`�%J�)]yxu��Ib��c�ct�N�P B!����^��ܧF�q��b�ݿ��}�ZC�:��p��(����G��Ш*5�ޔ�q�y��]$c�8M�ѥ׉*�����ݷ�s��Ԋ
�^\7�����bv.��@ĪX��<"Gn�$��H0`L{�Fx �&
$#�8�H�D�k#aa��ڏ;��Y��a�BsxI�2\��33"��� �j�	��hK*fƂ�1�J�ք؅ְІ�#0K����"'�*$�i�""c��C����B��iIñ�����"b�d\,�/1I��:G�ÁD���Ʌ���!�u1������i�aPA�v��I2\��5.�u�bA���%���Pt)����h��AM{�&"�8tj�^K/;�[�.�Y�k;�ݪ�P�]s��g s��Z�;l�9ܣk`^X����se��v60�2����
�3�h���9�l���m�s�-�P�s��m��;m��`c9���%��:Qjk���������@����OrH $� 	$�Hݙ��zM�I{�� {�@6rN��6�vZMڨ��$�.�}$�ޒ��݀	�S��O 1`ak�4M��d	vqxP(�؏0�.�[t�j�muLT�h��\kʛs52����lf�0Բ�70��`Ť�ͫ�[�p��l�V�#�5�jl]F6��f�k��gUƣ]�0&��fK-34vn���6ڒ��PhS����l�Pp�j�b݌� X��3vrU��b��7(�Zj�P�mʔ��ZJ--������,�..��h�f�Z65^Z1+6�� �V�ш#�1�\���mr�Y��w�p�Ѩ�ѣJ5���hh�ۮ6m�[[v/��I��lŶ�F�6HW�M� [6H�3�Wkibہv+�h��$��K�J#�j�`�)q��A,��zɃP�vv��!���w1&�Im��y�Q.뻻���f_uʲ0�ڋ}�H���*�g.�?}~��N��W��[�����f(L1{��͒`B(�F!d�F��6�K;;�,�f`��<5�J�='s`�v��x�YGl��褳wU����ٽ��I��uo������YG��=����ODq{I�8���Ү
>" ����~��]v{���-�v]����י�"�Kq�+��uU��]}�y�y�}W�]�T�:�g��a�uthx"�dN�P�ܓ���E�$x_���u�'p[�y��*ĭݔҞmX���U(���&Bn�D/�%ѠU�(� ��!AI��,n�{��s��;�}�����Y�:z!ն�B��S�.�J����'�\��V����ק�W2���S�u��1#d�.��)Ou��#�=�|8ov�a�yZ�o=�.�>�K��5b�ةu��X����{�_��nN�c}���C`��fu�F�Jɸ���b�'ZV�ے>��}�<D���ƛtP�Dªl#�H�jV�(�^o�C��rI%����v��A2�6-�\���їgiuJ81pS\�.l0lJ.a���MP�06��T �"��#6�,$5�ͅ�m+K�;��>�=�1E�nf�B��H�h����� ���UY��nLͰx���	�8.����w�����r���ކ[�Cd�)"�N
,��q��DeoHɎ�o]�%	ko���,I�"�Q.C���}���Q��J�k�$bXu@���y�v6�=}�H��bLZ$�R�>����ν�Ӳ�x��Ȍ�Iv	=��8p��Tԡ�Y3vyF��󞓷/9�8O-��`��r�s-a{���z��㛪{��>���f���\����έĸ�']�{���?t�-�;G�%m�>���^������c��F/v�/���[5�:3� �D�B1��&� )��6���n\�N[k��0�ᣠR�M�Մ#����쎴Z��*5�p�С痛[z��Z��U�KS�p���B�I����2����oإu�GT	�su�nW|=���U��.<{�l|sX�r��6]Zz��;=���������+��Җ^oQ�#�ƈ��ݍ����j����7������Ν��r�E��d�)��Uaww{���k�E�r9]��v��)��-nI�ҬN�u���u�q0���֓lD����v�h��Z)+Ф؁������i�1��]�c� ��?�ﺉ�x�T��(1��r���wpD��μ����=F6�Cd�8��Q'��Iy�.����ee�N`�f�T�I�r-����x� L����+y��;�zE�=��w}��7�N��e&��T�^R�|����?��˗3�w�������5,	R���鲜uxjZ���=v�w�6{�/ko�$T^��ؙ3L�B�=��ugבN*k�A�c5 [���%��e�$���������'0�P���,0�A-}�w�w���ڑ�5X�RE��bu�wm�B[Μvx_���Ԉ�z��͵���%R�nB=H�	�^�懑-nD��	Vg�i�t�s���a�[{��3=�T�Z75SBj����Ul��^����<½��w�굾�A�g�g�۫��㩆�gon���qce6�l�~� x^^��NnI;GG���m-�;��]1}�;�]n��>ޯV����hZ�[�ޘ�y�۽�,پ��\��1*����,&"b�E�޻��{<��}��'�NH���I���W�9��S�k``��%�5�X�v*]n�	ۼ%r��x'��9������O{J��I�ݓm�hb��Ш6�2)d�eI���$vt��K3vPRAv�w/{���S�oo�<���rK���yܷ�Q�ETl�lmM1v�k������ ���{o�}��s�~ႊ%θ�:]�͵l�4�3u� W�#U��q�ZL�u�n��@����%�n����ı]/"�f���]�;H&ѻw؍������ Ṏc���(��J�ܶ�P�j���������l[�lT,M4�U�onS��͍���Zf�1]?w>�:�����XU�W���)H������X�z�6V5��-s�Rv�"z���I�1!vv�e��݌��i��~�=�"��sw�7An\�̜w������?z����+�q����쫕���Ia�$�Pʿ��ܷ�b�nܑS�d�(���՛�gf������N��+"� �+=ҬW��ER �-%�*�	ZD�l.Kc��~�޼��|����v�z���	����_*�%�e[i�26���3%�I#a�}GMܸ=K��2��K����Qi˃1������ܧ�����cXB7\֬��4ҿ{ї�#$�i��U��q��;ݵ&�!�j��s�ooo�e��]��Q-J�ʥC/��Z�����)#8�zFLj�ٗ;1;�:9�L�Z�U˻��1sҋs�W�Ck8H��mVXx�6�Ynd�zG� .^��Vrt�Dq��6Yתh��TEJ�ѭ��O]Ƣ�R�/{���t�����Ӯ�]�s-�]x��9�_Oݥ��=i�P~�=�J2(��i�R�iD��2��@�iS���^�v-��ӷt��ऎ�\{2�'K��R;�s�$&�̠���R�|�UR�d��G�n����D��y;$����5V�w�� ��� ns��eH����uY��ں���5+,�.x԰$���/q�R��va�̧Q۪�1���H7����RL��,�}�  ���Y�OI�:�3XRS�����tX����N[�&���K�5| ;�w��&����똊�T�bX�S*�����?�T���j��эͳ�D�:�룪��JL]lJ�ɺ������#�v$#r�$�EI��-Qm�sHD�3��u�nwwoY5Ld�Z9VmZ�@�s|b�73���g�y�n�^�z�Oa�B��I�  @2[���e��Z��`�uP�7"�L<ڱY: ����V�����ʇw���Ȏ��e���י;�1k(��7�T�ݺ�\_����7y�_X��񍉅��'C]�9�9#��+Ѡ��, Ci7b1L���[�	y�׃8���[Gx���*2�'A �ɵ7�������ܨ��wYb�)�n�"��>��3��T��vU�0����yc51����p��Bt������e\�&e�*X��hb��:���x:�c�:b��J7s�BZ�q�vt���7q�T�Z둩�fԯD�Q�8�|�$��F�s��ҡ�37�m�fE0��Ă�l���F�6�yTP�r[w94�����U�b-�XM�4S,��w���%Ģz��g���CnV:��)b����kt[SD�n��ţ�lƅs]e�rs"�6����Ɩm5�׊��^6�f��M��}�nk	�����l�<"gk�����u�X�I�T�|��� �WW�i�V�v�m7p[5�c�]~�ߺ��Ǒ�U�zTk+��g��B�$��1l��%���6oO"��R=�&b�7lϺ���#�X<Ey��Cn���^������}u
H��;�Y��?{�m��{�?|.BC���Sua=�pW��o����_�o[�/N�xq]��r�UX���W�zV����r�鮍�� �չ��^�ml�Mz`S��7�u&�� =yB b��)��m15币1(_߿O�Ͻ��6}�w{�����������!��?�����:���-� ��D@��d�"��ǿ˂ j泑�"�UC$�U �'�Ȉ	�(hPG�V��:��B
/r((��T��7����3˚?�$AUD �ϻ>��������?�������.g�>m��X:?�g���K����=a�������?}�?�A�!�;������F}���o򇿣��3�Q���������Dl���N������D >��@!DI?1��������;Mf����3���X�?����~������g�" ����Q?��'/�w�u��6�p�?W�ρ��f���G������_�~���������y���4�;_���_�?����}v���y�f�DP�X  %{�A?�H .�V!Q!	Ea	 D 	�!HBF� 	d	$	�$�"�� �� ���� e`a dYB� B�IDd	 !	a	E@�@�!P�$�  �%R �!D�ʃ 	�@�%D�$XBD�!EdaA I�	A�$P�% �$F !XBA! YP� BP�%	RP%H�!%�X�R�R@��a	eEXT`BA�@�	DdH�P UX@�T�$T!@�VD �%P��  ��@�d�	@�I �XBA	@�@$�%U�`B�B �X@�<!%F@�dA�F  X@�	B $H�%�	D�%X@�@�F$$D$$P!	 ��	`%�	 ��	��	@��� ��
P)�@� �B���	��	V!P��	I@��aQ% Q!B@ �*2(�� ��(�(� �����*�*$���"+�(*J�J��*$�B�B��$���� � H
@ �*� *L*�f���<�?/�o�����}���_�d@D �?T�Kw�����`��������f���k������t�>���u�s��{����* �F������};�y���'��?�����7f��������+_���cߢ-�����?/������P��o�>��^��O�~�������?@D �:������㟻g��}7�v|���o��~�{��A�" _��3�m��;�s5�����;?>��|�_C���4u� 7�������y������gxD��}C�]j������?g@}��;~��ZC�.����볳i�iP -G�������������~�~�<4z~B���:?f���_~ϧ����������ۿ�����4���=9���ٝ~�������~d���ϡ�?��_�Q�{2��@���������~������_�~?��z��������������}>��W�?�C���������8�����c #�k������:����?]'�����۳����k�����~�����@����Z��м��?~'��s3�p���l]O�{�~��˃��}>��vq�����?A�PD ��~��C�}�<����������~��A�>�Ӯ?��=�v���z��O=��7�Y�v���~�?����~'��������d�Mf ?��~�A@����|��}��Ox                       ��ֶJ�Ü�^��(�          a;2�2�R� >         z#&�V������ ��S�       (�p�٠V�Њ2�	j��    ��b0q�y h� L�֢�F���AS�A�0m�l��N�%�%�2vu�F !`d�� ���y��s�������US>��**T��γ��*%�H�l` ��� H�� 1l�  �`@��= �}px����P� �j3� @ �B�!v �  �u� @ �(Q� ��f���5� ��DA!I &�UM`���B*= ��q@���ׂ��fP�E"�j��M�R�aI1���(*DT���8 y�0y�l4i	���J�J��"��"�CcT �Z@��<�S��UUI���2 k )�*�J�*�`��$�U*`�o�x�1=��):���UE�I�j(���(�tIID������U�2����|�[�"$�U ��� @ H�)@�Ң���(c
 �홈3NE��H{ SX)!*T�"@���5� * E鄀x       CT� ԥJ��  �� ʟ��R6�UDL�	�CCLS�*��UJA�     *����U&�M4�1h`��C$mOI�zh�yG���5%I@ h   ��_��}~�\KZ���N�\T�����TP �~s E<vpШ�y�aîyDh�D?J��}�hEPA�Q@0������O䠂 �+zDA/%2P�߿�uU���������,���G��C��@ë5� X�� !6�4C�\V��C�m�h��Vp���!ά8p55՚�� 58�rph�4&�f�	�a�p��l�C�S�98P��4:����@�� :�D톸@��!����6�A�M�8�A��h��!!��9��xւ��x\�x�M9�ּ �� 5�5�h� �MC�A9s�?@=4�N@4                           ��  j �7 � �  &�@ր�@��P  �4 � �����k�Ǥ�@'8|x	�R~�����GǴ�>���z@���Ƿ�Ƕ�ߎ}�>5������Vh��V  `|@�C�  
�h� �� p�� Xh�Շ��ÀNVx  ��A��  
� S&��zyY����  �Y�� Hw� �n��  k}�|zC��~=���zp c   `�� �v���wXh���  ᵀ �� ��6�  ��  /,�۫?�C����<~?ǉ������<x�=��� s��M5� PDM��}@5  ѭ �Z  $ �P  � �M@45  	    	؁� hZ�P Z��� F��MC@ j  x�d��BNM@�� 4 &��9 ����&��54C�5�hxx�9 F�$�55 �o� Mp�����f� 6�� %^�4B�����<�'*��h�
���� M�4�Ն�d�C[Y�A4�|f��ּCk	���7ɮ^#lᣓ�*�rp��7l�p�*��Mp����9� U� X  T` V  X  U� X  U� X  z�  *� k  
�  *� k  
�  $  5  	  �  $  $���G��VhO�<M��x�ޚ��<��湠 �P9��������rHr'k���@���� ���9ANN�sG!ɩ9�h{rC�� ms�� MCY����� 	58��9�4  I��kG=5�5� sG	�ƼO�CG5�G��y�� �H                  1�   0`  �  `  �  `  �  `  �  `  �    1�   1�   1�   1�   1� ��c�P ��O` ���m���]g����׫!�`d4��@< z� �m� c �� �� 	�0  c  0  c  0  c  0  ά` �  *� �  *� �  *� �  =V  ` �c  ` V  ` V  ` V  ` V  ` Q� X  U� X  U� X  U� X  U� �  Y` �� X  U� X  U� X  +    1� 0  `  �  s�Ϗ�|���'����z�}�=��C@d ��@ � x ���� d��O d8 �  +  m�4 6��#l�p�@��� ���#�> a� �ٮ������>��@s�yf�@�@��h4��>ì�p�X�@ d  V@ d M�l� ���8�<kƵ�� �l���;��   1�   1� ՟o���m�� ��C�A�`���,==�c�=T�x����Y���` V v�@m`��c  0  c  0  �1� 0  c ��X h��k  
� X  U� X  U�  U� X  U� X  U� X  U� �  +  ,��٠ d  V@ f�l��@ 4� �  �   0  c  0  c  0 {�&�ğ��� �d�}�C�yg�h}�~FO�C�?<��x'�V{|��{~��� ?����fsZ�30L�3��ј�MkBfiOy xy@���В�Cy i�ka���4Z�1�y��2R��)JR��*��)JR��)JR��(�iJR�I�I�I�I�(w�\m��۽����OF3B�p��J���D\]<�v���F���,�Snj�*z�JVl��:�"��ERO\*N�W�X��T�L�������8�]�К!�D�2�H��p�t��Li	l���]"�<<bYP���ܔ��"�١�� ua�u�����Z�33K��Z�}ff<f�rVYw�N䬌ĝ�'�A�غ�E�rO�.�4�m��k\~u�0��JB���)JR���Y��ݩ��k,�A�y�B��yJ_$�O,�['|�,�y�rI0������5�@��%#A�ݸzu��2���A��j0�,d��G��B>X�e�S"� �"(�*j!:��C=�36�nc�n>�7+q���������iJR��)JR�JR��)JR��)JRP4�)JR��)JR��4�)JR��'���o�u�Xg�}�<o�q/�t<l�f'���xZ�HR�E�o�����JR���	����<;��R�I(Q6�	*R��9*Q��=&"n�-]�&�*��\��R�5��]���i�V�2��l7nC,���� ��(�с��j\�t�NVF���>YhZ�'y��{�	��f`��&���30L�3�0J��30L�3�0Mf	��f`��&f)�c�����1�c�������������K**��A�{���DN�����e1�׺w^�)��b��1C,OUU-�sND�2w��1X��ݼ4��*��@��� �w��8��禷�q�˟Ւ�!�He�d�Y	��C,��$2��C,�^��/�Y�h�NZ�F�o��Ϭ�/��e���~�[�(IT�SEE"�P��S�	৥E;��."�TçM)�&.�����Z���,EKҪ�*`�)S���5T�-��E�S�YQB�vI)�!3D;K�H_ i�<�o#d<�b�(�YOoqV��S,$��L��C�X�������<Iw���>fY,�/>����ܘd
��1�2"�j� �w�!�(q�<��dvjh�!�g���i�!��q�<˔2"a��X�ww���f��P�R���k[�;7n#f�v��Z���^�/[�^��2C,��j�DjթujS�V��Z����������#���ѽi2�B�)�A
 �����ַ35���kw,}3Z�̓� ` 4�  *� �m`�6� 4X h�� 4ma�ǀ+  �� �  �  h  H  H  {@�  H ������ D���<x�  H  z@ @ @ @ �        �                    H  j            � � � L�     �  H �� �� �  � �  0  c  0  c  0  c  0  c  0  c  �  � �  ,� �ma��C�  ����@6�P� CkP�5ٷ���Muf�@��g	�jk�!��  `  �  `  ��|C\u� ��� j���!�h�CZDZ4 ��h4@@PԐ� �P@k@ s�9 ��  ֦�M_9�c�����$Z�9�5�S&� ��Z4Z  'Nk�9 ���'4hC\�sF��G&�rMr�k����h��r&����59�rh&�8��p����h���D�5'	�h��k�Ѯx5��x�9��4rs��4s\'!��5ɯ\<�85��4�]� r��u����oXUQ��G������u�����}a)P�Bw!��'����Y	BP���7	�J��>ΰL��(J���J��`�%	Bu	��%	hJR��(M�P���:��%	f	��%	�M�P���p�w������Q�!(J��(J��(H��(J�J��)��R���M�d̄�(MBP�&��n��J!)"r�]��:���(JY�P��� �)8F���;J�%	BP�%"j��`���)v�%	HfBP�&�4%	����p5b�y	�x'!(NBr����!)J��5	Bn��'P���(J��2��%	A�قP���'P��y	��'�`�Br�N�7	Bj�L���%"d%	BP�%	��+�J��(J��(J��(J��(JQ!��t0�DJ"*."�wٞ�#L�haPæ,C���Qe�l�(�����T����:`Hr	*�`� C��L@��%�^�=v�/'O�Y���"�{�N^�S�w��p���hd���F�c	֍��x�cOe�!ϩ������nBX��_�R9H��D4'I%sJ�)(���MG��CR�4M*�XP�YE]�9��F'e�� ��br0�3�5Ó�g��|<��'}^0z)�)`�N&'B�ml)�I[B�.{��ek�VVX8�U���r�jU3�S;3�;�m����L�Ү>4�du��Ј�T��<�Ȗ%�pO)U�j���w�L�W��mX�MD*S 䒞w)��+�l������FZ@��Fsa���on�N��o�q���yw��A9�B)?�����)S��$	�o��9q�Ӿ==����Dil�̝�,�f�ahe���ҴT�&|��
��P�R����9	F�L����9	@a�`��� �F`�2B�5��i���p2�i۸w�R��F�w�7��t�����H�}�I	'��:)�V��p�x9M�ֱQ<:� �g��0�2h�2�	2L��2)��� ޤ=�r'�ɱЂ�e"�Yz6�,nU@ h���)�s��|Ǿ���S�,�)Y	BP� nBP��	BP�Bu���H������:��(J�JR��N�2��&Brp����	�MBw	�%	Bd%	Jr!2�J�Jp��	BP���(J��;��J$4�n��7�!(MBR�J��+ �Q���(MBP�%	BP�%�!(J��5"nR�C!5	Hj� 7	BP�������{ߜ�3����3033�	$����Vfs30������	������	���{�� 733���znπ���E����30��q�ݞ��  [�      ��    ���   ��      n��s30�2�=�&ffff`&fn�aE �> [�����;��330332I-�
(�� �n Q@8����������L�����$�(�� �n Uz�3��s>�n Q@9&�s3033330     $�      ���  ��         �wv         �� �       {� ���L����{�fffff`�H-�
W������f`&ffff`l�333���333033330+3,=�>����	����D���L���f`333303$����p{33������H��pX ���3������L���w�����L���30n�(�� �n Q@8�,�7[�0���{3333033331$�@2IO��$�L��$�-�
(����|Q@9�> [�������	�����������nffs30��U� -�
(=�vL��f`733��f`&ffff`&ffff`�g� � (������E�w�`&ffff`&ffff`&ffff`#9���� ���� �fI;
(�$�        {ސ  fff      ��     |*�w`     g�� -�      wv=�d�]ߜ;&ə��ܜ�{����L����˻� �� ?ff`3��߀   2T�0        n��  �     ��     ���   �݀       Q@��     ff`&fffffI%[���`| > [�Pn�����L���{��33����C����	������	�����$�> [�PL�����y߮��ݑ!7�)b'�.tM�9z5U��̲�(��8/9�G�_A��D�(�<�v��%D���=������Ce�y���R,�e�C�	-�2�WZ�����C��9���6�}��}�&��Άmb��N�A7���l^G2�.�m۾���0C�̒$�ݩ#H�zi���<XINؔ]�m�}�o��߾U3�h
�����i���=��㪨������ﾷ���Aٴ�f���Y&��U,�wk���_�{��]��ܫ��8��{����=�Ro�\;��p����9��UV+�s���Ĵ�s���B��s�:e�s�t� ��߸�*f�
̒6�mɲ:��CsZI:�8IT���ݐҌ%$�����  Fr���v�b�>�i��j�c��/m�F,X���`Z�F��s��Av�c�u`s����mݒ�����aUU J�����U��l��M����;ޭ��˕[b��y�ޖY�nLS��w����/{l�ƿ���� >9Tgy�/��E���9�0�;n�d��ΣE6�>�ݷ�_9J��,9����s��lI$�[[Xŋ���{��b�6ǝ{�A"EVd�%�(�t�AH��m%�v}�M�9�V1mc������1��*��t�)�kwa��0`������1�]� ��o���vյ�{��t�"������v���*����UW���d @C!�UWf�EUL�����|�U@U C9\�����
w��>�N�-�����N�}������Ӫ��]������ww�{�]�w���߿ ]݂�� �� {ސ��Wd}�/t����Iy���m����/$MUf��ܻ�����U��p �U̟H��ͽ�UI��� *��� ધ8?o�� s��~��||��Ϲ�۾����p_7eW� ��ԾU]�7���4.���߮�>�y�$��}U�� �*�۾d���[;'�$��w�w��\� 
�w��{�p����K��f��d���=v���*��v���>�s�ήs�]��9���͓3~ߴ ����9�9�UW�RUS�;�.φ�����_� �� ��I|R��y����*G>���  ���ګ_��m�˷��|�6�l�N�}���@.��
� UUw������wO��*� ;��{��s�*�����w��J塥�m�� :a�y�{:��$�2|J�����%�Ψcm�l�fN���*�뷧���}  {�s�q��@UK����kv��Ty�[޽�{:��m�z$���������w�9��T��g9���f��ǽm�޻�{�{y
�����Uw�B���_.�|}ʓ໹&fv�bg�� U_s��^��*��I9� $�̯��q��6���;S��E�������5���*�����������2Iݽp[m[o2IU���}�������n�M�IB_rN��ge��I&ۙwG�v�飹��-M�Um�vh����Э2�9�[/��x��&I#m�ۄ��7�s0s�=���0��n��w��T��}~��ﵟ^a�y�����ʫ���Nng��   f� ��Uwv�w�@�>�U=�ɻ�=w�����o� ����l�*�77`�����}�ϣt�'�$�*�I&�mk�E�jM�v�agr��E[:ƚ�Rkl�wN�.��âd��C����q�>��띭��u\�7o2]�k g39�����}��s�INv��_9��URv}9��wqٙ��\���:��<ꪕ�#n�ά�,؄��a����r��we��z�����j�m�T������E$����B���}�sj���$����H��Us�{ޒI�U[h�w�J�������uU߹y�s�����   ]��������|�9���{����|gd���z� |+��=�w������� 﫽�@ 7���ez�=�� =�ڪ����$��|�s�s�	$���9��� ˻����   uK|$��N���>�͗q]� ��T�� ��� =�O�� �]�I!UuWUAwK��$�'8  UW8 *�� I�T��*�������� �������;��$�U]����p �ܒK�� qwvU�Z��&�6��{�o��}�)w_��zAϸ.��TI��IwvUP��$�T��>    ps����� ���g��l�T�{��z_sk�z   ڪڪ ���w�e~�~��Cݳm6�D���.]��iۻ���2L������� ����(���������[U�-�V�Uv�@�^}`]�U�| �����R��ϔ}C�����o��������s���w` �� {����Gw�}�f��� � ͒  |    U7w`   ��  `/9�{յU@�m�mW���ww`|���]��%���Um�UQ������g`m1y��s��VԳ(l%,�
��Q)<L(�.^��w���^ �?{���#��f?�I�������m׃���{��=�t#��<�}�23�w�Il{��=����c�����Sض=���%�ֶ^�e۹w��{;���wN���ǹ,Ǳ�ga��>�|�Ǯ^˸��ff7��6]Ǳ�c��e�}�j=���w��{�{G˶<�}ǵ���;�j=�콏��ձ�{�{�[Ǳ��c��%��}$O��>���c�^�����{��l[D�bN�#���%��z�_c�^���;�j=�n^������=�l�����˻���{Ǳ�z)��"��l����ҽ������wa'3v���w��r_.�{/�t��ovw]�;y��l�kuL��J��-���w`         �݀	$� �O{�         ��         ��      >   �z@         ��          �݀   'wz��z=�G����z=�G��vI��� �  ��߀   2I        ��         ��         {�         ��         ��        wv      w`    Ugy+��>j�N��=g�R�}[�l�-���8��+X��oo�^+}o�s��̸�e��wjt��UQ3�Nˤz�_"{�ke�t��;�z<qX��YՁYۄ�c��J���6��S[��Ma�f��U���r��:1:<�k��3��+=�&�����z���>���<���N��y�ﱓ�|��tH/�z��Y����[�W�1��o�H�^����t����U^�YW���m����:F�3%������4�N��^�,�9���½g���p����)oU9��"��[��6Gqb�7�p�.ٝ0mjCk/s.Z+���z��ܑ��u��z�z�N�n�W�����ݺS&�Qe:-ɖ���:�����:5nT��Xko�����6I��os33/Ǳ�k���˳�+4U̵׽���l�i^�f����lz��3��O=�^Wz�;�PVs��fndW{p��.�ly�r�=[�ww�c�ջ��=�c���n�ޝP���=��UD��Q�yrt����V]lZ�ug�Y�{\�w^k�{%�{6+�l����>��^n�e�r�w����ɷy�L�ocٱlym���V�{V�Ώ��z������귳33.��K�u�M)���큥7���]��T�����VN��s7�~��^����z=�c&�3�d���ڂ�"��;X-+��9���r��_4��Ⱥ�W(���X�w�2���Q�5lUU-��n�Iff��ŊխW�e���9�{:,�[1+��6���Ι��n�C5�]�X�j�%d�o&�d^�6ӻ.�N�q�$��+Vݻ���I>���9��޸�S*���N�;1�z�r�g���K�n�y��m��L���6�qNV�uW�`��.[��=�c��=��O�b�s�*�3��y�[����0C�̒$�ݩ#H�zi��}�}�~�C�L���&r^}�ވ��4��y�Ǟ����TP@Pg`���[�����Q3�p����v�슪�(,��݅��-ʾ����v�^r�w���y�s������}~��@P��s�L�A{΁oi=��d�zG7��z��|��s�p���i%�!�JI	$��e���}ʾ���!������-�ŏ�����1�c�s���Ar�ݎp�(.�,r�qw��[wd���;:��UU@���|um*� �Sl�����h�r�Vب��t���f[���������;���F��[UUbݗ�����vRы�kS0�;n�d��ΣE6�>���/��M������o6$�s�8�c/�}�۠m�@�u�׳��2D�ĔK:N �ZM��Ѻ:G�=�l>|s��>��o99�ϟ|uJ���](�`���s�LʪTj�b%m[X��O���m��@@��UJ�UP�UP�쪠 �*�Cl���2�Z
����oUTUP3����J�yyЧp[�����b��~��H�����~���Wl����@!w|���*�����n�z ���� s������~ 9����߇���{�>�
���s�_2Vgo�Z�����^��n�Ps�Z9��W9�.� 	��̒K�U;�W��9R9��8  ��'�p>I9�s�r�3v��[�MR�̼��f��/2H�2�$E$�NI$�D��ސF�nId��w����U~����{��wd
�=�_��
���ݵ�U ^s���{�Ψ	��RD�7T�J䑷���SẔ�{��W.�>r���U�.�=%����s� UW���W�6
��J�<�w|���V�+Tf�m��T��s[�a;wi$�}�Iw���S�C�9Xz	(ZF^��d��}�Ĺ�sI�Ĕ%�r��*Λ�l��l n�j�s�p$���s� UW��z�eP�-{��rs� Us�������Ͼ�*�	��w��U U_��Ͻ����ހ  ;'z��&g]�ޯ{wwә��L���,0 ��`TP^o��AUN�E�pT�@���*$ ���� }@VQڂCB���qP8��"x
��UO< �NmbA���tt����G�״�:^�]���@|PP�b���*���E��H	�(�P�P< � _==w�����hi�'WO���)�<@����Q�z@�0��0�U�@�I���8 ������x�ox��:q;�<�;z�{v�'���)`�Bt�}�p�;q���*v��v���xo{l1����A�N*h;��6��y�K{��:T����Z���ң�t��6�����Й�M�X��� z �/O��E�3� �(`�J������HH��NXm�ڏ������y�ݱ��<KCۀ#�;���/h}� I(�H�/���I��] 
��v������18iֺS��ӈ����ç�!*x�=�z�q�^��	��	����P��:=T{S�;��Ov�^�;W�4mN�:��0⏎�%Q�8$ ����Z`D���@���
���������'��{�](�����7�q`_�@��z��z�i{�(�"������������
(�~`�(%	�Q�A�T�AJ!&��(J���%�PDP��K<���_��G�Uj������.s�ª����ـ{$� {� 	&� {�n����<{v�8,
�{�ٞ�{�v@q��� �n��� m�w���o7���]�� I �@$�{�ܺ�s�U�\�}^�HB���P*�/ev]^-,��䄕Y�z�;����7�
�E0�I��"NfĒ$�=���ۻ�D�7e�=�w���u4Z2�f�1�Y��8�B�I&�n�F�Q�rG�n[��2�v�I�Rt��渕o)���m=��G�5$ǌ�˥g-ٲ��e�M�1)C�?��sg�4�G�t��v2��w]c�LH��m7�w��q��7xc�J=�ZN�a�a�*e��Tp�hݤ�uz<�%$����2�6�7F�6JJ�gg���1��&�{��4�b���?b��;���ND�Vm��f�UC�pr�O�W+�9u�tt {f����p���$ $� 	$�I �;�_ܝ�i�e�������5�-B�%�>T��`�[k��m�7!��.�w�ݟ��Ǚ�����IU׽G��$���QvI32$I�ؒD�G�X��C�wr��Wm[ӷ|�&*+��5:=7�Q"ۦ�$���z;�1*�S�-�U��IQ�@y�ڳV$�J$�yu:Jּ󯞛 ��� `�~>��t*|_��؛��qq7֑4��1S��QG���ݽ�Wa�1$&���lf]d����Z��I�J�k<�Cq��5.�l�*�I��i�l���!�����U��^L�xf4�a��V��\����[ߪ���
B���^�^�T;�۠p�/�q����z����|]w���G�6���Xk���v��"x����Y�1L�0��>�nd�]��8�ad��BL��c3.FE���F8c�E��6X�36FQ��e�e��6Fx����b��b��
	�9��aَ�q}/x�Ϫ�3�Z̾�2��ś�;5, 0,��'AG�3��]2p8=aл$�fH�`�@��u�}{�𳭓��)4j1��$�Nl�M��#�1�lĘ'$�0!1�I(!��C$Ac%������Dc��l,,XD�x���T�(xL�QLS��q�d�@a��IfgI�l��,,l��lY6�A���7B���..<�	B�\��t|��K%������.i�	
sV���#*��fc#� ���2r22�����O��I6NT�c9�)8�Y��2\�,5��Daf�5f�	�	&(N&��o@x��L�d)JJ22	����������
2Ǒ�``L@dIADHL�ĥ$AII@dd��N*�y/�~��H�B��*d�&Xͦ�#0* ���0#V1j1�����6FNXYVX�ce��ab���X�bŋ�b�q��ܯ���XXXY�f��c�c3���8�A	�:
���{/ވو$�0cx `����$��
fA��-Q.z]>>='J>*�� z���"z x������ >���tz((�(lP��^���O �=G�<N�P߈���z���x��T����C�S`���� �
�=A;@�=UW���/�=��/;3�5�tm	Ǡ�����<���N�UB}ES�T��:wێ>�уDݡ�
�$�i,���^���� =�dc�%������J�B�N�1���==S�	�&Y��ه���"��f�`�	�CcǛǽ��ww.�v��a���=�R �tlN�0 ����[3&aFM��Օ0� �6���r�H�ԑ;Tҁ���"h���܄M�,c������~SblNǴ��HQ�==��͙���5Da[����;ww3g��5���p�9a�ZD��}c���;Bfa�r�̚��j�f��]#���u��=è��4�bK�+�!Պ�ժ4�<�YysD��iB�`�NIP�<���43��o�y�22*�ZH�Ȧ��`�R�Q䝝�(y��0�I��kEthڀ�ە�6�a?�n��>Xc���2]�)����%7��r`AX�T�vm�+�E�	�{��򱦐_n���E1��d� M��}�{9�ܐ��$�{w[o��]C�rf��q�M��۳�\�P�kM��v@t�#y�n��\���p��7���/����3�w%�$�WS9�sL�'*L���M�©�8�;�DX�6��f=$�R��`�a�9����mkЉ:0��^u!u�܄,���2�	����.ـ@�+�<˽3Bu %�gxp���@Ó�*5pÆ�ю�%P���{�=����˼��5��GfY30j|�ff7"a(pށލ� "Sް�5�!��b��;T߯fk7�I"�5������T� ��6�8s\$9�-"f<:8 i�@�������S��&f6���.��u�W<Рl�`��w��Q���
�ݣJ���`�����4
��������\�DKݝ�G�*��0E7�B&��}�&��14`�H�o4xt�$+�R�f���6j0YD��&o#�r�F�{�[0�AXI>�)�0�f��U3S��8��B6�Q�0Vd[�NyY�Z�����> �/J���f��IY�T�f���]����os�wsvcKX��vfr�7,뛻Ѵ��n�]���)ӸA��Ȫ�S�z��w����P�Ȭ��� 3��y�{wu���_<��):b�A�nHoFK�b�'\���$��TCMG<1�@�|q��;D�LB����BB��bM�j1NЪ/*�c30x�`��n=��ܝ�kX�8�G�D�#�h��kP�@+ūw�9b8����U�h�����AE��MN��N�>X��D��aʆ��J�P�D�r���swP����� ��=C���f�U'gb-��Wo��5wTL�:� ҇j�PU���'��=By��U8�i\�Tvi;���M9�׻-�t*�,��I����]���ϟ_�s�M��+=�Bu�N�G�4�E~�j����n�u�;=8P�Z@��T�&i���5N��X�3�6n��(�ঝ�k�m�q*�};
�e �}�VP�^��b�r�:�@���N�����D���,"L�*�̚'߳6j��J!�z4R\5�P1H=-f�4	�Bj�RH��2�4���q�$���V@i�˭�2\�L[y�]�S��0�T	�0���Cg����g��u�u��}�:rZj��ݼb��5S밂��D�='���őd;�+U�z���;?+¾���ҫJEn�7v�U��h�Q1�j�PJb��k�~��v2�F�g-�\�N�QG��C�V\�\z�5�.��%^���k3��"tL�5�L1:�0�� �E�v8x����b��{����s�}�~����m.�v���}|q��z�qjI-"�Vɍb�sTڹf��ÇЉ&5�w���y�Z�2�Q��޽��zyţOV�� +�x��f����M�7��2�L�la�#Ҥr�H�f��gF���몠��#��s�L������/�k%�2F���D�<�3 �m�GE��r�)zf���_}�h��(��id�2����^l�^K�ӷ�v���M�%��K �YySD��H���ۻ}�O�J'j�p��$�o�xr�c3!�m�U�I1fX�S9�^ݷt፵�*\��CJ4�V��z�0y�@�1K3���� �]�N���(�yu-�t|jH�7���_|�x�(!�����DzO9$�庸>i�{��z.]��Exffr��fM*׻վ���画��9ͫ�
����0H�iB�Fd�m���׼����]��6�w�nw����t������md��{0� ���f��y�wr����v�/)�߾�;5ETNXc}�r� �$H��%1�i����kw�e��I;x�^$�����(��Xa�P�~�v�*D�ֺ��h#�����]D?���yI(	�A��O�`墑�e�DP⺨غ�]�fդ;����h|�c�_������%v�S�U@N� �,P\� h1A���+�*�/ue1F�6�_� ���� Fa�]$����"�ul�Q5�%����9V��3������"ٙ��ܝ��Ю����Ƹ^{h�O@���#�&�+�Gbͪ�*�3,bv�ˊ�0A��&�Q��� #q�I|��Nx���$��}�Vn�)�fe�׽��Ի�m=�Y��#ϯjm����<9�ݗ���ފ��1�!���0�y]udh��3 �>A4�sQS����%BSQ��w��w ��"�y��P��"ܼY3臨w,}��8���5{wFşY�1f��_?uߎO\ֲ���0����4�3�
��F\d���=�o��t���4���l�ʕO"�2�	�#�)X9��,���{r�ZN҂��-�t�ϑ�9��b?��U���.�����-��IaC�M(5�QKi.���8Z��|~}�A�@�2��	��,��yӷw1{b��C�Iǧ��xB�Z8)�}8��O��0ѩ��)qd`qY�]$��:��{�c�2���z<�6w�ZJ%T���9�/33��ۮ���\�*�����e'hܝӪ����q��R�X��|�~����v��d0Tv�[tE0�j�ėv�乚��]d�����H��Cc�f�Mg��I��1&0c�~���K���7*u>��xw�G��&jԖ�e�G:�3
�4vG��-w�=�5��=�ލ66-y�4����5�t�ʣ�(��a��D�0��xw�9g�sqȔ�����IE7��RCUF��fa��آ���\:�ݱ�XC�E���,TbP�瓶��ne��m�F*���%���`� ��e��ة�H�Z1	�d¦r�>+����(ᆭ��J!�R.U<�D�P�W$��[�� y�.c=��ln���s'9�e���%��w=~P�A2��-�r�ѻZ�f&a�#og�!�
sQ�"(v��k�MS�#�1�Ɇx�1�S:�Z����fM�;���y�����nwwi�7�&7�*W\̷����2ʳJ�U#>D4�[�D�乫���b���y�i�ޜ:)]:-{LN�SI����ˤ�i� ��nP��)��������B&ܚN:�|�h��#�>oVV�n�]Vڃ^.����069B<���%��
�����S�6�ۚ��E&�H���-G�*�A��\�33��)�*�bb�I���e��-�0�NG1yU��ۻ���&ݢܘ�V��"�x�-;�n(m8u�QB����˱�H/�BU���2Vte��ń�q�`�vw��(e{� }��:DҁJ����]�2R^ܙ�|�`a�0�C�EC�xM�k���%����Z�����3V_�x�P'��k�=�UL�Z6{s�g=�P gP_}��9�wbF�BJ�kw�	9�zǛ������M�S6f�y��f��n��ۃ���7L�{���=�ٝ��+M�%*ÁP����T
0�tE��!�ŗݗww|��E����	���
A���:L��;m$Ae�4��sT���ﰷ|D�x�J�1��	- �NP��G���^�\4#:�Ҥ��;���WP޽������UD��`�^UQB�"c`K<���{�r�u��ÓKT���I�R&v�p���d�e����p��"���4fa������F� s�ql|{�e�_��V(�"��xv �s����=�2[[��(s�LcM`_;("�Lg�E&`��$����fe��K����D�Ў���5���L�p�%	B���	BP%P�"�%
�*C�(4(�$�����i��� ��6�#I�L$���e�%�`�IĔ RĦ\J�3X��v���%<6�!(J���(J��(J��E(W!(MBP�&BP��J�����ϹϾ�?����� 4?{��I3������$��7w�303$���>7wvgnH I I �7vn���I$��� �H�$�r�7wa&��(��l�̓�  �{$
� e��˃�� �H '��`;��I�E]/Wy��+*����������]�*�36�R\�٥$�yXP7O�]�c*��$�]�t<�:�K�us�3C�Ns��7�>�q�q7}�U*�� �*�>���,QBzl^�V|�s�8���R��7�ݸ0�E^��������ٞ�sy˻�ək�õ\˪�:W,˗��^W+:
F�sܗ;�ݎZxC"�w���]4��ZS�4��*��
�؎��ЬeL˫\���cd��$�1d}p�Uʮ�#i$��ݾ�������
�f��l�[�wO���c��L	����y{ҫ�=�̒�w�ޟc�p�|����f�3���f�.s�.s���nös3y_[�]}�q�}W�=�~ ���d�I  7w` �ڕ*��;�  �d�$�*���-�};u�+Gu3�r��J���Q�5<�P�*&����Ŭޖ��]ַ���43�kf�5�l�m��b�\�G�l��R,�vsuGd�����[t�+0���#3kJ\iN���t�Uئ2��2O%�7C̣���W8���|�Ns��7�>�q�q7}�U*�� �2�	z/t���yw�U����ו��Qm�xM^��f\�*�u�/7_L͓e�{׽w��s�r�ח8*v!��eCn�N
�����&��ʿ1 pdAd��b�<8� k���;1,�zAm�&��TI��1�#�u;3�Z����V�Բ��v�q��J\ɫ����e��{�I����T�&Ǉ���P�W�D	� �A:� B!� X��$b�B��@Nq�pI4A�8A�p�!H7w�=�AC��"�r�8�o�!�z��p陙�^�{`�A &�tl���b����r�0����q!�@@�)�L���/��ۻ��:�p������=# z�(:���XvB!> C��8� k��b	%�P!�L�����w�<�Ö���b�!�L��j�`�H�:!�Dά�A�o8`�&fs-�c��S���}�z��JuN�a"�@�9.��'(BD=@a�@僦C�~���3�c�4�8�iG�?nowO�=+����P���mA][4!�w���H�qў��x@�Bd��7ad����6w�Tƌh�P���@����Š C�V3�`�z�$�@AD8@ra4Kү5�k�ך�V�&�؆�s!l"3j�3!7�y����l�0�����&m��à���]���UUZJ����(!I���C�F�9d�0j�xnd�!� �a��GT��^��\�g{�/8����kA�=� h��y�f�^��1�!��7ðp���%T�s�,;-��I8�$��If{2�쑣K��o�©3.��wEՠ��s�g;����F�tb}�s�{w���ޝ�SWH�j�%A��h]U՚,n��e�3����=J�S���O^<��4f�������&fB;2�� ��3!�a�!�tA��� n`��C0tx��f�aǗ�)i��$:$a���~vC�hf�3)8:C9;%35y�[�����\m�3`����A�kC)0�|#�0��������� C  C��!yy^گ\�����|���y'P�!0��-���C�~�ta�!~@a	�Xk�	�5{���y�i��t25��`�s���:#D!�D'0�fa�����q����d��r��x<!�P&\��J�Nh�	~�Ph��VPl��b�R�H�j�W\�˪c�[ �6ZN3���#�>"�h�9Ճ��=��f@H�G#Dv@���3�A�@r����3���>�W�4�<���P����F�+�ua�7�`�#��k47��wǬ���њe) `�k�����"z�X�Q0r������l�!�BC��~a�l��g��}�Op����� �xp�����S04B�z0٬@��d���M����w�ϐ���3�٘�v��EvѴ��}�{�1�}�"�ŧ:��1�D�Xn�m*�:�F㾯����e�z~�'�v+���N�Sws�F;�1��tnnT6ro~|>�/PB��7!�gf�d!��>A�^��L�F�=C@�1&jL������N`ށ�a2�8�DJ<"�`� �d1�F��!�jCx��Eȑ���z7=�����ԯ��
%�8y��FB|���̰`��zF��A���C4@���&���,�鈳Y���H� ��wP!�9��e�ry+� �8��ϝ�#�A	�L�;׏S0��`�NP�r |��f��tA�/py�) ]V��7��: ��h��We�3X���������뻻�<x��Al�q�0��y `�iA�z�(�	�	Ơ52��9Ð�!�`o9������7	A�b3	��C����+o��c���ƺpge1H!�����k�4��x�va9�ޏ��!�Qȁ㎆qtF�'Rò�0���xD��8�1A"�0nD"Y[�q��wq)ޖh���h�òJ0�;�0���,�Q�Äu��NA��=�����J4C�<3o����荗8q�JC����A�>�0�xM+�;�כ�A��(9 �-��x8�Cw�#��C'eݍ��	+Y��I��2\�1l�JUr��f0�N\J%Zf͛��I$��l�1mⵏ{�t�x��[S�0o'mf�P��zF�+�u�a��9�`���P�A�:��>	�׎�aL���q���]܅�Q0n�Ӈf��da
F�_%tkv��2����� �^�{{���pŠ��� �3�
z[է�݃��؄Q9�0ެ��ž��+�?o� ��n�$�w��s���&s��S.�X=��F�k9�3T�+�yޖ`<h��dq�� ��=O������ʘv�t��n��O�CU�s8�e�B�,$ҜH�p,��>����9�Q��/6ȌQb���ns݂)�M��ri) #�+/ʉw��4��V
�OP�U�WvD�
�MrL��I����*|���ͱda#��2����=+��ݙ��=ީ�p�3�E��Y�"�#"iHTA';,eW$�-�7�\�0��c$26���}���W��U��üf���&�")�&�!Ӓ�Q���ضr�۰�bf,[�c{-�s;z�nnI�9�QI������O�w�,C��S��v�b�b����>���k;gg��|1�}�2�Y� ��a�M�z���9X�'DYD��A�7���v�}ٙ�y	��x���܌�~�$Ƙ:K�'��30I30�Y�ΏL���i�{xtC�b;S��c
�kIc �Y�3��b��G�v��/:�j��y˂:h��m,1�9p"�f���]�x� r�oOoF����܂���X"
�7�W�#F%�9F9@�8��s�3��w���VQb��I;�� ���s���&������(�����وta~;:]�,L���/}��E��qʮ���w���3c*aL>$��xFP� ��O�G-�� ���� =N� �v��7���̕��28���a��N"lNs�JH�$↠��e=�9��vkl�J��1��ǝ�׳H�p>��X3Y�뼨�W�g>������x�g��~ݺ�=���b��D�͗&����{Ϗzw^�&.3�Ee؝b��V�~B0��WH]��eIT��I�a���H7TB�59�O"��E�O��(@E�?3��f.��s4f"�f�AY�ADa���辮����im�J��s�a�ʵAqC3IG��W-�rH�*�}��ظws�;q6!Ip9�8O���'�<|�o0+�DMWGBN�Xbc	��H�lr��'�,� r�A~�L+7��US��� �1SD%��0���AZ�x��4�D�s௷���]�D�|H�9� /�EY�3��Z������|�IEEI%\��[�S��wx��E���r�@;���.,q���V���ߕ�"�J��k����8ag�	�a���� ��=�����_�Ι=���(�	R�e����$��9�zX��m�@�Jfa�r�=fg/ܜ-� 4a0ۻ��S���ͬ��J˻WM�Y�\�7t�Z$j��\��mb�!Y��h�Tˢ�%�+�KR.���I�*w��{&��祂����$W���N��?f�d�[�W�`/����თ� ��������|�o:W��"h��x�;+h��k�rE���H�OJN����˻�ц�-���s7�)8����&�fbH�qFc3&� �=��Y�w�x�f��^��Jķn��d���I�xD���q��EQ��[C��9���d�#��*���r�]~��Ql�8���o��{����5"�Hz ���<X슸 ���R9b��00�8p/T)�_tvdW02G��pD� �d�yl�Q����Y�339�� �W,��)�a�@	��D]u�I(��P(��ʰq6�Z�'DYD��A�f	$��}�)'6����������t+�"[ �;T���0A4���|"q9n8�sw�����ܛ�6�H�	8�rܫR_��#�02ˏK�T�Ȅ�u\���$!%URI!M>�=^�ߝ���n�&>���Q�����s5l���]��/��̭Z�Z%�}0>{��$�y�wrˎK��]����}�ʎ��!����4jA�ĚQ�9c�O�Rk0�Ab��@�3k�a�u^��gbD8�%�\���PЅ��<�$�����泹~e>pTK�Uvl�΋3f�#���u�+��o�h��V��x��O���fX^Q'lK�w�H�`l��]M�\#,vF�y�H!����I4�6�/��e�ӐH�K��%@�H�٪���yY���<W��5�w��94��}�Od� r�T�iC�w낋,f=Y�n}���ݢ���8����{7�)��Dj��@M(O��P�@���q��بT.㬢r-d ��^�J|ga�P��3V�" �����T����1l����"�~����P�zX�@�;�w��
M��Ͻ�2��C��5D��|I~Xa$3�r$�m[���T�cy���ݹ��ù�i�����e]ݣo0L��kbǵ�o���wq���$7:�f��$�Y7V��l�\�-F�y���Ϙ����ġ߼�����"tG�)��d��A{ĘRNe��3$C��8�2����!�P���Ҧ�Q�����
��Iif;��z2�.zH/�<P�)�{�B(]�,�B�?3U|�����G����.\϶�c�8?�4	��=�8��
G$r�9Z�EZxh.���m2�U�V�N�:�m�3�[�!�
p����0�͝�nS���9`!�OyO/W*�����xO�"Qc�Q�9xn��a��
J0=D�A۝��먮�Q/���d!�l�S����rxE�-�N3�҉)��q�gLΈP���]�iDېO3�1˂�v��t`�qbs�+#Hw�#ii �ĘQ�>,��(��'���}%�j���"����{'34"U�Z�%��yǤ�	�X��ff0��3
��q�A��2�C�S!:�Z�RϽ��Ii/�w�3f+����vfi�/�_]
�V��$�RI��b�f���)�Gn�0oH8p��j���E �t�	0��|��&ý{�t'V�#�O�so�>{��c�$�W�Đ ��E%v�1�,B1�*�k̔x����d̻�@���l`���1����)�}]�lB��sv���z=���^N]g���w���,���i"6Р��[��RҩL���D��-��w{r��!�9�P@g��
I��Z�)�$�Ri�:z�<����G2�4B�=I��=I�8���'�,�ҷ*���fZ�}S1�0]�@�����	��$BK�v�*ӋS�J��OK�T��ۙ�7'�rr�#�b����+�^�X�2�ƐC)Ǉ��S�sq.��>ԋ0�϶�N�ĎZ�q��=�,��2�\m�x��3�3 i��p��^�IG�rn+�8���? ����ǻ	�A�<B �����B�9��'=�����A6�i_@���Kf�a̄�H��,:A��('�"�H��;Q�hJv������SP�&BR��!:g�hh��|ֈ%g|�����u��1o8����"�eنȜ=��|���su�^g�k���\9��<3����}�@UTW�6 �H> �z@2I0 {ޓ���.�����-�_W���30I$��� �n��� ���� ]݁��� d� I �@$�{������|�9��}��nʵ\咫���7FأU[�$�lI���C�R�M��bk�I�i�(��ӥ���U\UP��beUP�{�9:D�rF����s��v�{����~˗[� �ڴl*g:���;�L}��]`���]��ϠZ��g=Zz�d���n3v�A�ҳ�N���Zf	̚�Uٻ1��&e=0]q�1�òoe@��vqں�SggpDM�mW{.�v]�q3�g9-�ȷve��l����%�	=l��H�(���� ��i�F�����[Y�u�M礪u9i&6��5�i}��9�K��fћoѵb�����L����>��F�	��6 ��>��.��H I$ I �@=�H��ݴ`VR.֎ʁq���+X��7x�i˷�r��������ShHb�S]߯~�{�9�]mn���ؒ&;͂�n�X)��,v�������ݽ:Zh�UU�U	�6&UUT37�v$��nܢe3��$���DD�ki�}�ڮ��]�$�����i'Г��	���MM+��Ң/�`vT@� ���$��4Ц |d�
Ș(B��
x�Tt��:4�a�30��Ь�R����Un�s1�wj�{[��rh�NlT���]������*_��l,:$�`���ޟ��Ȧ�J�Xs&M�ݫ�B8od�ь��7y�z=�mG��|�˝��S����]|ш��4(��	*o9�h�q+94��y�������|��d�9E4$s��	Ļ*��f��$�=Iu��t-���	���A;�"�(�`� ܃0�G�<P�!�e30�F�{�^��.�9k�W����E!�D�DqC�&��v뺧�B�}c C�`��p9NǠ�&�))��H5L�F�����.��31l�#�A�W$A$�*���r��6�,��r٦m�޿v��ϙ�TZsP�I̴��`r���tag+�砂iS<��=�Vw�hG�$�S}à���("���y$I� t�ʵ%ɾ$�ܿIQSoq$;��J���� �;q X��P�I⋁ᙙ���p�S���/'+Oi�$I�zYէ�݃���ƣXa�07��d���"RviԄ*iif`I�i���ۻ2f��wy�iv�n𭏢�F�Æ��ynÍ��׷���N�t*����A��wT�E&�n�������Rd��2��	�@�˂.Ӽ�H��q7�H�I����4�}��߇�"e ����Ƀ��lM���x���0{[#���g������9\M����Cq&���{��,X�����c����{ww��x<㷜�`�SM��94���ǅ�@���L�L^6�|��b*A콸(�����S��2O�I�� ���*A�T� ��P�E�@�de
��D����8�VemO�/��Om{c�*G\���!�T;TA';"p�$�'�D�X��� ��Y������`�;Ye2�����%tP���Dg�<r�]�m��D@k�R@�:�H�e�l�H�$»�VFz�uUU[��H� �r���PE�6&�3�O�N'1��fp�>���3'{���$�&��Tm��96��p������V��eN!�5���Lm̚�n76��xs�{��=מ'��Q�CJ4�	3������]V|P�ۉ"L(�JܫRXI�I�=,�Y���O�=��%���<�qZ"��3X���T����.,q�s�H�	f��FA�����U稻7ެӯ4u���� � ��0X����zH-����M�7t^N�F�A���ZN8�Τ��C�0!C4m��?M�:�f��뜵+��G�(�ILS���t`��G)�d�q�5�?�<F�ҋd!�$ҲG��H0�k�L	
�p�%�{����ں�B<��W4V
"�@������{�:�z�wx�q0+`�vt�m�=

 �V�$�>&8���8/u���0c������Ѧ��t��LzW�&�`�<v�0v��fr޵�p陙��H}��q�P쉨(ff��'��qva����h�'��$�"&H&&a��`�`� `�&b!�"&"h��" �E%&H �XBV���"a`  ^��]���m$������9�����cA�[2�{�����Y�yvv�X������c2�������n��}����p%�I�ȧT�lY�x$u�y�:-'��)y��Q>��n�p*'����㿮"x��i���"*ռ�K�UF���^�b\wy��u�F/C��"tE�9�U� /~$q�r�m�2\�%
����cLK��A�Pz*�3�_�	�|P ����{g�z2y��EId�����R^Y�\P���D�Q�[��^|l�.��AJs|�����8��A0*z^��:El���{��p�&8��=���P�ͅn�����^��몪�;§q���G^0��,���<�腆,a�=+�=���ڂ�a/�9{$�2s��dp��d2�/��/c@�k$�]�*1S�k5�%ąt�K�M�{������b�e����f}.ȋ�riI�!ox�u��Hu�9E4%���I�f��ɡ�_�w^��Ve\�E��)���ibҲ����F_DO�q�1�ͨ��Km*at�K��CN�E�4���̗��&�N�y������I��K�/F���S��hܤU��6�[�)��9E�9�d`^W��ʣX��ĸ��*��%K�{����(��Hx��Q�z�q.��B,ElOCjD��q�\��R���%�Ij�U�ۗwkO�d������#<� �V�A.$[ҩ��;�Y=���ms-$Ki#�94���x�
I̴�$��4�q.)�ur�zfJ�i6��nr�K<�Z)9N8�'�"M(�ގ�����kP�R�j$fa��4��_IP����Y�[P�jr�յ��픒SO
�G����EQ�9c�N��&C�K�=ZxiY�u��eu��{�J��KA9n8MY%�F�AfQ%�/��]K�w���m��Mάuĵ�D�P@MS�?u�I���ܐ!����g��w�����$�iRS��8�I;��z�,���ܼ&�#}5���k�$7rn��vH{��f�]��Q�t=ң�>���=Ѣ>-��t�9~%�Gd!�I�|>��[U��xf�Ffs����� �S�.;s��M6';׏30��b8ruY �d�Q�>,a�qb�BEMɈ`�aC� �<�� �fe��,�$���q�p�z�X�@��e��\O��W.���<�������x����t��N�I�dUA��=zyT�.�{���A���V!�\S����o�j��5em�
�u�1��ڕ+�h����	�DU�y �h��Gy��-�]�u��3������<����{J4���I$��("Ĝ�f>���{�0����*g�,��NS� ��$I�@�[�jK�|x��
dҌq*C��Q-"is����ƱՀM)~$ �k���ؖO��=$�ܚJݔ�۹h�>��\�]�N�u��[9,g	���+��s;x�ܺoisz����v��oM�������08��
�`[di�V��$�(���sg%=�ͪ�ff�p��M�0���"�;�K��r�M��|�]aj�n	�d�p������(s�0���k��2����A*�� S��͘t���ѯ��r�"!��I��ь1�DP���g{g����O<4�DVc�K�
���������c��R@?�~RK�z����b�]�ْa���PA:��%���޼��L��q�8�Vm���,��dv:�8�08žH��|͹����;�T�����n�5['��)�6��G;"j'����s��5�c�_��������\c�����a\��$W��/L���1�V��|��{W#����-'-� )����l}:�����u����<�9��f`�p�kww*J�/�C����}b�cch�4��-�����߻�>��d�勨�*y�q4�*Gy�e��^���^�Ovm]33F�*����˿�6V�ҽ��%'0sXbr�"
"`�\Y��N; lJ�����7��N��@����9n8�V�M'(�GK�RP�]r8�e�.��J����޴b"�
n���-�@�9����.,q��o�z_2���8+	�W�f-T����:���q�O�$���$����>�w��i�>$���"�;�K��zI�yԎ���(���ܮ�و�"�vt�f
uz>��$s���
�8����H�����ʘS�7�QM���Cq'��P[3%N��� �6d��r�}�9���+ׂ��!��n���9T��	5�R��8�`���o>i�Lh��<cA�\[�RN%�Tm+ i��d���yNEc�ɣ��t��+}ͫ�DxrM sr�zO��&)\� ��y��j!��!$K�%��y]��Đ��w�Sen]
rL�7�ZQ1H]�W�Y�S��n$���DΗ����r|}���s(
̓��f��r���*��댚���jڪ�,B9��NTA'��6��Ҩ2+�5�Γ"�IY��g�)�K��,� (���_+%�l���e�s��	��	q"ޕH�e��I�BrܚRC|��|��Nn-��"��mNש�I�H`�\W��Ns�JZ!G�I�'�9�z��D�q"l^��OY�nU�.q%Ź}E0�"�S՛3��(]'il�b��ȕ���ė�8��
�`_yo���S�I�rqv����:�f�H�98_�I|�t���^q�޾���=	8��N�wRwx,�����&[L�2�݅"�A>U���-H�qTk31�6�y��$s\��
�<K��F^�:L��%��f'��RK���Д5�a]��W��0P�f����� (l���������[3�s��DB���m���.i�6�ߤ�Uf&���{�K�Ug��W��đ��E��杯z�*�9oX�ǯ]�:˻��-�U�SM��8�R�^�(�@�e/^{�g��<���Y����..������f��jd��3���nP�9G��X�0�yg����$�['�\X�p[38R�Vե?����!2��Qws����Z~N3�<H쉨 ���D��c�=��;�\�{s��"��k\��Y;D��2Mi���儖P���H*ռ�K��TE�L��
��������L�����)���S03P����Dt��#�N�S��~�r�W=AD��TbNlJZ!G�I�~P&��d�3}��nNp�m&�	C'�0A�^)2|�%��=g�ĉ$�x{;i#WMs����a��2�����rv0PL�A�[k�a�u^5�g<�w9&8�8�+��Q��f�9�Ai����N��> hMk_� �$W�S���I�D��rh���D�B|���I�6��J�	���C�%I6{18�3QF��BS��2���k#*!L\�u����kKٛ���OWfӆlME�Z׻�{��ho}�$�70v�� ���[�0�����X�ݙ3�@$� I$$��=�x�d���{� �HNrsܩ0d�z�} �I�&a'�@��ww���UO*C�� �@��$�L�̒H�k>��gԦ�G�g[�j���"!���V��y��u:�Q&՛͡yzV��*��ޢI���U��Ъ}�h1�[�(؝�	.��Թ\d�OJ��uL���*���˪���H����M��Y�:�t�n攞��T��Dۖ�X��wҎf���}R#.RW{ww:���^~x3M���(���G铉F�<���=�o�>s����ۇq�υ�-uȸ�X�*�B�.�2�8���`�j�M"6I#l��]�uG*�_m@�	6����{}�o�{̒�[N*��:ʵ����.�`j�;l�8.s�v�Y�g9�fk��9]}^�� {}��� ���n��&�J��� �@$� zo6�5��)c�5�o����:�+QD���VZ�e�*j+�S6U�� ��]�!Pv��vˉ��j�lÝU3@0��>���{h�rND<���#�;n���I�f�h^^���ʭ<����z���flt*�u�uV��6'n�K���(i�n�L5���uV@�a�{�F�-��(�vC[S�ꤳ.�oG;�����z�݋�Z�˿ <E]�q� E4��8�	11�4���O���0)�ǋ�w��}�}����\$�U��r[8��w=&9�����V���o������3�뛻���[��m�S�}9�헹��_��xV�D;�J�}1 f�+����Io��U�QE4Zߧ����uz�_��)��*�=px�f�L0`��#��2.%���2�^����AŶ�i[�Ff=��A��,[�A.$+,���1a�2�i�y{s�#Dz���`F�h���Pp������%��~��:����������-�`&�f�:S�e/L(%��S��wX�@�X㛐G��O�#�z^]��_|Q.+q�\ ���P���&��HND�2 ��#��T�i,�� ��ĉ@:,zW#��(�ĵ������]��(s����sŘe�<�9�J�H%��0mFe3#���-�P�^�M-��V��Ƚ�$��=0��"J}��(o����˧�?����zNS� ޤ�M({邆�ͨh&/J�[��y3.���J�wٙ�m�˳Ӟr넚���e��˔����+�[32Őr�I�|ֻ�5�f�9����L���nt�_Ì���.�I���;2��}+��2��^)���l�0/e�/�$a�&��Gam"�ʮz���uO�}13����N�a⌁�r\҂`^�/F`�/�d�ﯖR�'\�R�X�q�q�G���"��(�v�N�G����=��S��ʮ�x�5:�>��d�"�ܹ����AD�9�&�'����먮ef�1�����:L�W�I�A�6�iO���U�8�Ddj�D
֣`���`v���M'8c��ǈw��i�P$_�0� |Y�Q�0$07g('�+m<3��l{�۵���Р�s�yN ��C�Y30�39����*�8V�zy���>*��	R���յ���GL���Dx���ߋN��x�H��a�rĉq"�*䂝��^%����|�$C�a����yfyz�ov�Vmm�eݫ)&�ic�`�ui��Z7g.��̤�+1��j�tP��E{��f�B�mS�T�J��L�r-z�q���E��\�UT�~�c��O&#�&��L	��Gy�[����������{r���9�RCb�iD9��d�$�ܞ&|�I�NQ������<���x��Y�9O*�I��C� �MFɚ������1�-RD�^���q�im"��%C:~%�O�^������˻�G�4����^Q�^�\��	(���Vx7�q�H�HG�ꓽ0G��e�H�|�>�=�^�zI,���T����A�")��'�C�K���JB=�ǽ���"�^$�V��"��2�B�<�{��F�٪�m�~j0�Ȋ��O�˰EE�QT�����v�ü#�)yZ$��)�}���R�l'��s
	s�0��$�0Ã��_���27}�L}�%۸�owx^�j���&���۶�B��1���aR��۪�I&�$��{�����{��_j�z��)?jcs(B$�oT:����J��g�osݗuŜ��%B��d�"Q��A���'�}yo�J�u���}�"��Ҝ�V��섪�$W'��a��/��L�kJ+�]��T�R'_U�i�����b�~���kj��c/y�wHS�X*�G>��IՔ��o����˶���F5�V�<�Ro]�]Z��|Lʗ��b�e�C����J_���ȋ}SI���>$tP���������=d�h��U����)+�y1�z�j3*�w]N�G!�n��AYWUACO��~4XӺ��.K���1gMQD��'�������m`��[��dv�$˩��؜�ؓ���ٝ�ͬ�]���;z��|D>���ӖMջ�<��3�����>�{�Ubڜ.�f}I.�Ŀ'CaƓ� ���$9����eLn�wn�0��"|���*,G�RvK�qۮE�=�Oz��M���j��c�a�.R�|���w�!�x�i]��_�"��z�׸�y���EF{�P��[~�{�޿:=��W[WV�-�%Iˈ8��4�3;�e�=���ʲ�^����#
f�_D�;��8rʨ��"�O�6;�'����Ń�*��+t�i�i;yWp�S�
���ꪫ�fc�1C�S�D�E
��1�"i[�+%��1^Ϸ�ou�gj�_�g�M�ɫP"��*�p���"g�{�L���\_����q��b,D|HG��Q��K�����K��Ù��3�(�<V���ۑQya��V2쫓��m��TE6SuK�����}��o��V�����¥���Ć�d�]�K���Q���0�Zq
�?�_����"Z�+�$���9ޞ�q���������D���I"9Գ�?Y!VfT�d��㶲�]o�]�!ᴬ�лE8��Q�^a��Ә�x���p�O b��
˿U��i��yvdFn��W]�^�j��"�=���L|���7�Nb�jj�umD�7��}bW��B�z!�־�s�3O�O�<o��OF��35�i�፶ލ�m!a�;/�,5�^�Sz*��7���ݽTOj�wن�z�H�VG�噚R���|L��W�tl�t�{e>��c5M�y���b���2y�o0e������V6����e4�r���[�d�W&i#G����:�EJ��^M�۝ٍ_�ӟ��9k��<t��sZ��7�1t���Dݔa�<D��ӱTK�sLR���f�#=����i����E�1y�ڿTC�O�vR�����g|�t�x�T(�!zȵqX���6j���/e(M}�rEX��%�.�^�z�����	�cG�t����Fl+�vz���9g���2�m�cG`�"��O�LS��x_�e�u�ύ��V
�r&��k����������Ѷq�)$q��Aw
���Z�QǙ��1��<v]9P=�w�����u�#]��yz��	�R����h[���+�U�Py��u��z%�����h��65$;����ݍ���n���݄��<��Y'>�~�N�;��F�঎����of�Đ�ɻ��j�#�}G�7�� �<��%�z�K�}v��Sl_x������U[����:��'d�U�Ej�5�%S�[�'��7���S7괚c9<�sU}� ����nԪ�,��<��,��F�F���"M�]��Ʈ]�=wwT��n�=o����eЮ�}�~���0�U��=6��HF��1�{ř]&]�y֫[��-��Z%]��b�z�U�،Ü͵o4��}��z�F�gF#'��%�כ���}�}���yl��î�Y��$��&jb���Iq��Z�����;���uj�&U1+��"��Y�P���礌6ri+uD�2�7.F挝�ܭ��=�0nي�7=�e�rg�i̚��ٹr74d��7"���iQ'kªX�wPV��۞���n�ޱ�}����az`���(��5P�ީ����{���w<��s���]b�L���U���ީ�DU>�f���̧����w��U� �μ�l��̌V����c�*qq� ��*���0ݗS�U�y�G$����<�:� !������,����]�H�����������^R�gJ�j��cPy���~c�3(W'H>#�ڒ��e���rR���0M�ʙ���+1n]'�Y�S:B�3�&ĳ#b�������v�����N6�=U۔s3ي��V�s�=��|r�SWeա�L�(�g]���I��1L>��{U[7~ߦ��¨�-\|�8���'�m�L��P�ej���l�}bv��nǖ�QR����
�	�eO-w̦�A.�v<����[�'��ym4�`���Q�����	jx#���ɁULJ�v��l�0Ԕ	x�u�$�^�	�&G�<vr���SU��v ��!�Oz7��U3�|� �yo��/�ڪo^��U��m��ǻ�2�b9;GNN�o33 xxF�qY��w�͙�s�;��M|�q�a���>���k�L���"�V��̺/�򖻑la�v�֓HMZ�fb6yMN���˾�NB���.�����"����%DG�7�.��RHSQ
�G��T�[)6v=ը��M��{�0�F�8�!߰KA⇡��uh]1��m���|M'	p	�3AkDh��)��d�\����&��: �����.���d%BY0;��^6<u���6�����o�`�11d��F�� 1�$����������,�$�Lι��{�W hJEh0��L��"��o{���}����� wg�633��� {ސ vI �����}�b�����+��UҬ]�ޑ����E7wa3306rH ��3.�`� ��L�ܪ� ;= �H I I �}���w\oxs��T�w�_ٓ�\X�i����Ecu&ȋ��N��K�.��h!l�;��k
I�Uq}���	4ەUJ���ꪸ��s�X5N�o�������{gyuv��m&zX�b�e�I�
.����Unl5���Jfbsu^��D�]�6N��3+y$�mv����7f��G�1��5g#}ܹ��z�D�����	:v�� ���Zjv�<����܇kV\�Y8�f�e��:.�͐L�s�|�mU����
:�qH��.�EmP�N��H�B�ɝ%��S��|6P��wq&6��3�ҁ�2�&�����]���m�|���g�l I.���$�I  I$ $�w�A����������V��8���D��#���Z��k�f�C:�X��y�3��ĩ���m4��ݔV7S�D]V��+;d���5��y}aI<��/���a&�r��CZ�UT�w9i%��I����Q�3��6�a�E3�=5���n�<��v�A�8S�%�\!�BL��ԏs݄����]L�jY� ���a�&�0���cX��ӂ��)ڎ�4U����[�{̾�%��3������փ�8�ź4t�PRF�;y�CP���Pj%]���^w�96��	fSx�w����\��"�!�����v��9�Up��h fH����31 ��4�t�E*�~ލ�_2���$7k�ի5lc�oQ[�B-v���s{�m=BGH���%�ioE0�ϝSi=��͵X�gf#/��j���G*�E�����^�����k��U�a�$��< ~�o*���`���T� |�������\�}7��zcaSb�0�I@���%ـa�j��a�c�0.�dZ�x��Ֆ�1J|_�{gL��C�+}�.Ɛ�b{UE0-}+«z$�{Z�V�柣6��gqYZО�PN�$ WN���2�-�Y�g,FZ��߅��i�O;bQ\I˛	�f茄�m|�3�Ɂ2`��R���y�9�<��}$�Ifv�'��K�2d{�$�ApҼ��)d�ɩ)e���HI$���l���NfP�����a�`K;#a'y�0��Ǫ~�;i���C���8�r}�,����:�~�Y��b�\LR���n�p���/RMl7�{��]牃��^�-��Jz�fagA�z��%@����R�G�]?<�ET���V� ����1�=ս��]��Dئ8�ܾ�����U�Hβ}�UV����'���0y;��^lU�%q)܃iF���#�z������g�����BOg���'&
�ŮL
��b������n\�W��o����	zx�u�e�dT�b^�����*�����3Ku��� ��}�h��j��ML$��׹��d���4ܚJ͉#Mʽ���b��f�{�������F��K�1��o\��E�{�������'x��� uj�����5�<W�� f��);����CC���|��;�,�r���+�e�}�O*��Vw��{u5�o��i���qeO*0�< Dҷr<$� ׼TE�])w�x�	*�Myk��i�5Wxr,/�쟫O\��ߝ�s/����ۥ�qlYK����+�&8������MGO�j.��`��x��U'Yu�z�y\:7U�<x�-S2Ɵ!�3aR�{	��]�0��d��Q,�]�E�a\�6-��\G�+}��y/�M;t��O���eI��rE>��s�d�V{�̸�tdWuTc�U�}���*N��b�٭�Q(s���Lw�ì�6s�0�,���Ȳ���z�_`����g9 誤{oll����j�Wj�b[#mS�h�t��a1h�%��}��7�`�Ryf+<H���/�cZ��s��rݯ����F�.i�3��F��Bϯ���y��[Xx�(�|v��>�,���~�*R6��[���ʖ�j��/PsXM�|Q�Q�ɉw�n�=«z%;�����0cG�N���A��=�O���x`'0�t�jP3�M��d���Ṗ�z��AP��!\�ħQ��	�eTM�u�ޅ�^�3n���=Q�@�{G �[��YZ�EQF�x������U<G��Rm"�u�q흾���py��Z�D�u�T��O�vT+����oO>=0*!��L�: YV*4��:ȵV�ӑ��M��07����귞�Kͣ�Z��Y���J�2��rjӢJ��U d���yn��8 �#��o�Fˉ�����O��s�٪��ɯ{Q���>^�ʱ�}��
@ 5����u3i�8�t��"U����X$�^ERP��'Ž�yG/W*�����i9eج�:�������f��>�V5o��4��x��(�y���hf3��UgD�#����p3�}}\����'�|�TާòVǈ��J�)�,�ffY��m��R[>{�]=�t������SG-栊������xa~��Oݝ?=���0e2_,o
t�I�~V�\�
w�t�;s},�A:�TڪnY�-�_��s�w�{_�v�(V���Yաq)Ւ�e�p�*�k��ܝ�N�Ժ4r�nAu�R�Oer�kn`��~�Ϸ�U_�o���ݓ���/�>ؤ��k���;N$Oi};E�΀�$F�"�ޘ��x��ᳺ�<   )�EG���݀�<�����S���ғx���E�׶����ffLs��r�b]��cp�.��D�v�x�y���{�.�B0��t=�3��^x�S�mŦ{Ԭ���ʠ�TǠ�^#�z��5�,���V�B��W�r��fc^q봎l���tWP������D:��UG��uHP�G���^��}����oR�!��+���U<M���Tާ�N%�U�Gl<;�9ƞ�"]a3nW������7��. ����7�]�UU>�B�j
V'�T�^���j�ݻ~�җ?�W�tf�j5��kFφ��3~�5�ܬ@�$���PY�b$��W�>u�^ѝ�7ͳM�qY�)�j��^�o�Գ0�̰�����.�_\��˽ݑ��� W�[���{�������c�J�u��+uU7�zf`�Tk��[Q�ʞY~�Ѷ�f,����N�p�=�Ey�i5��1Sp�E�{wݻ���x�����`XH��t��i��3�[k���wXZa�a��.}��M��]�  w�Jܪ��U�go#/�3�A��*�_��.��D�t�x�T)�S^��i�;W-D���"�{�����v��\�֝�3�]ºC�$��I�b���{�+1k�T�kvǸ�-�e�͇F�lM�ݟS3>��׸�JbOƓ��. fƐ��|\���Q��ۻ���_���Tߓ�'Lz��ib��;��[O}����w�3f'|�0;�vfq�(ܬ��YT�����ӆ��]u��&�{k}��w�ｖ��6sv��m�_6�xf\�D�v_q�(�Ф7��8{�l�D��]Wކ����V�A���;�_ON�U1,�DEҹl�����m��`��
��@�oUs���]׵UT�omkC}�i!஝��}v�������_�z�\�SLw�Tڀj�<���WM��31���bΟ��ﰼ�fj�����4��њ4l�_g���w5�uUU��Ip
��(pf`�Sm ͱT[�q1J}}���U�yV��FX�[��p3x�.��%�<Gw/��+K�.DJN�8�T'#�#�t^�ET������g�cz䜴��-)�o�i�z{�UU]�Z�ۓ�*�B���HQR��`��H�g�Í��˿t~�����eݫd��{����)d�#��d�����q�n�c6p�E�L�!�E{��d��SA�%I��%���;$58�&���r�n0G���}����}�����mU'��ᘩ�,P�&pXXj�{z��CB��d���o�m\���{
���Rq.�Iv�Jɸ�z�}S��^�9Q��3��n ��(��[R�С��[mׅq���=�05B#d��q��Yo���뻻���V�����I�Mr��S?����^�̬RGk6��1��B�0�ՁBS�$()���^̜A�Q3�7�^ܪ���7`�]�PC+u��bu�-�)�l-S�Q\�X-�*���8*�Z9W���3sk�>���i��"�`m����� ,�)�C���`�_��_lə�[�z_sK�l�w�N-�ݕ�;���{�v�f���u9��`�I �ɻ���!z���7gY�f*}d�jژä��]X�-�i^F�w���9j�K��ҝ��1ޒ\B��W��.�����34�D�;ee��|��l�V�f^M�kp=��:�g��Ra��\V�̽bN�x���2rnK˕�Lf{��]���\�oSn��"ͭ#s�冤�Y\i%��)a��}�&P�����vX�J�\��7LҔr�`�PF����U��ʠ�F33�;x�I'}����J�u�!��-���Ϲ�[��S�6=�?��UPwe,���eݝ%��#V�a�N,#]�U;�º����V#d�$�@�b`�A�8�9�k�7�O�H]
2��4+��Dۆ��\-�f��Ɏ�o4�� (���P��L!04RuQ!,��oj��fffb��ޟI$�˻� ��/wv�fa�l���݉�I��~�� I$ �F��{��d�I7w` �d�6rs�T��I"d���E>I$	>� �H �yR� oeH Iffa$��Sn�ˬ���3?��v�̫�IKd�i"fC�k��f��8�XA���hS�҉���Z^a��Zi3�۠�P6����_2��{���I�ܣ/2M�31&�m�$�������Ho(U�ʐ�Rn�(���5�����N�Iw�Z���U��M^ɡ&��Z�Ǧ�{�+���a���r�:�A�p�e�E^�j\�.�dPř�pf��v�"�;�f%x���L��RR\I*�{UG��.�����Ng�1���}�ѺhKY�{{M�f�p��RS-RG{{o���ngH�I6��PW�0膵��j�m����G9�dlfg9�iB�i�Z��v ��w�@�� wv ��)�]��H 2I �@�ʑ���(-��֬��]Ga��āe��ᏚS.�	����	���QqMQ���ف�lS]�UZ�ŌͻXM�t�m6�&��g�I��������B[w�N�����;�(��I5���%��0N��	�oj�]U�+��Ld���2�$ݮ�WUf�C7K���&�=��F��t	5�&a���K;c�;��fm�t�Nmk E%��`� &=�@�L:Xp�Sa�	�e(z�� w-�4�c�UE��0�mɤ��{Y�qMST{37�]��3i��R{��o���M]��4�Q�bl]'�粚=������py����W��v�/]��y��@�0�]�H��|)�y��,��6"4pfbf���I6��>�.�������gwJr����B���]�j/շ����[�>C�(IO�.y��4��hB�0,�s���z���}�I�ZoQz�T�SFn��Ii�ְ���Nz^���6�~����dY}Rv?9$~f`5������{��l�j��k�dM$���R���6�U6�T��L����Ջ��S��{�
������!:�b�]�3�U�6x�w4�u��� �e���(�A��Qj}氝��U7_� �6�K*h���T�uWfQ�əw�/�v�e�ovGF�
�ZZ5&\��m�KuB��&�lR������X7i��V�"6��l��j����U��:vFI�bK4 }�̮���o�'s�m�z���3N���H��a��p��Dz���{B�_fSʻ��l��4��b�;���b�W�mx./����xYw��i432ח�N�����h�w��0*��d��E�e1��yD;��#�-|&-S�j�"�0�x�⟚��#7v�6�	�.���I߉�1׋ޭ�컺��j���.������%��-(a�˴����gH]'���Iq�Р����S.���4"� �+��H�R�y�#���"~;{���}UR�@�vkeO}I'��f�F�}4����R	H��k���Ա�ff+H�[���Ef�`��Q���6�"I�J�鹋��cW����q�DX1�7nL5�'t��I������}�0�{�N7�Q��s>[ZCB��qw��n�yF ^(���_�A��蔴_��"�O}�[i��g���nvP�/�ߏA�{0���|9�s��Qڰ� a��۞{��q�99v�t�-�&��A�RC3K���6�|C��j`��*���Ҧ��]��IEq$W+qe������H\*���2��)����}�ݻ�K�]v"
��^�a���v��mU
_� 3\����|Ğ�j�դEلP���,�<���C�K�T_G9pD/Q\fKS�JN�S$��3����_2���R9�+��f2���l�o�j�0
�Y�g�.�Ϫ���~�ĕ���vs4�*nM�;��Q�E�IK�S�f��U��wy�-sk�$'rn��{+��7rǫ�ڍ��a�d�=���m�T�x'UP+�lR�:�9��7�+�9��"��T��{�6�F�y�Z��}Ioe)@�N�x���rrb��s���f��ǋ������J.芩~%0���0�&;l�^#M���2�w��uLR�S3���_{���\�{�����u�*��}��|Rޚ|/Ԭ�~����In]M/p�*� �<�o@X ���[�a��SNߣ=�~����v	���Rc��-���ҹi3�u>�BN���]TA:�.I1V��G���+ܜ�t32�$/��L\��W��S>lX�(���g��_� �6ۓI[����ʆI2�N��ε�w>�vqO-�vk���,7���]�RI�Jv^�����9�Yܻ���8���1cȫ��,��eyX��7�ͪ�!��h��Q<..�^"���|[�~Cdg-s��&�B.a�"]^���r��6+̢�%Ju�ƪ�+�ؤ$x70`���'�*��$ISډ�rH�,K�Y�=�ȚI>ߊ��/W*&����?�)9�}����Z/sjЫ��t��V\T��[���y��^�8�Ԑ��W�v̞����/4�w4�s��H> �t%>j�Z���E�h�&�z��S��?\�!�*�Rz�f?p�����@򮓄S��SvQ������vc������B�(�#̣�.�f�u%���6���x��h�~2jK:�ͱ�����KQ��ʩ��vim��)�ISD�-�]B7�%�7d�:�m��  `o���t]��"���Q�m�C�XG�x*�D��8����I%2�E����I���V3 �j�U-�g�<u̽�����/Iv��[UB��J��.���]ݻ�oe>EU��NUv�N0E��ð��.�[���X���w�ҴX�AqG�D�{����׹^Mړ�;��4�gRh?����ދ��^��$p70`Y��V>��]���Og��8}��Nꨐ��o� 3x�CG���p�|�Y��b�Z��
�e�
z/�U���g/C��}^�7��擉n�IkHKH�wT�F0ל!�$ q2�=�z�w6*��~��f���M��uNI������J�d��.�m�*��/�)�D�k~E��n����)5F�5�l��y7u�9U��J� |�}]��������+- ���C�栍��ؘ�ىwZ����ռ�������^h�+" �` �=u]
�!�V�N��M�����*hbA��uϽ�2���ߦ��E�D_��ʦ�B�v\[���*D��0��,Y�<(��v�R�"��wSΨ����U�ꨤ�-:�8,�ks���n�����Nsg(���.��j�z���O�ɥ���ͪ��~]!��A�=����}��]��D�}�^���u0�U@�o�JW��yw[ď	��Ȳ�W�r��
,�	H^�]ݎ��!%jIn���wt�Vwdݹ �0İby���-ĄJ���7y%WCo2-�}wdݷ��^�����399��r몜���?jؚI>�2'����I��^J���n�N�V�X�ɁU<�G���L�=p�g��Q֊��01����xL��1�dŻ����{wv�U}d|��)G-栍�Ȕ=�<��B�z���Pe����o���9 �+`�����+���xP�
fj��%I^Sr=>�g��R^A��	X�ܦ������d�cB��U�I�HN�O��&7�[����z�i�5A�sDAOO�M'�$�(�C����S�Ě�30�MIP9��?���U߆c���鬩���y�_E���&��<+�M;�Ҩ�k�ߦ�.#�=_�g��ݵ[��;��i�4��+�e�s�%�L[7����z�l�y��UK�����ty֖����7o�*b����[��� a�`fC ��mwwe�w��#�`df�7����R����YZc�őN�3ʉ��\=
��:��9��`�lJ�PamO�~���3���]M#ȕ�̉�{6���f�k�BO
{BصQ���o�E ]j#ޛZCB��x���w��P��N�K����a��#�4�	x�.��[�1��V;�4��u�ҾȪ��J"Xg�k�O��	���|�����]N�����>������"g�>�� � ���fjǬ|�(w��U���f�����A��p��o���)��z���/7ed7yE��n�o�{ݚ�%�;��陙�u٘/3xl����L���d���g]����=�#qv'���z��l>��:��R,�&��}A0M;Sް�d*���y��f7ї���ݜ�{�"Uf�>	��,�݄O�G�]�F��:f�xbL(0w��Ȼ�i�ޢHw�𒚱OQ�]�N�);�^$�f���{g�͝�]9�҆3
�1�#7�NbN�9k���rpp�ޥ�JKH�B�а�����'�Q�.v���9P��G5��,��[��T�ϩ-z�B��N�i>�����vf,׈�Z[վ���}0�3'�.�QwDR���0^���a�l���:꜖f�������o������]�W�K���6)$RO��E
g�@o7��]���@5_��@��� "� ����O6��l�*�$tc��ߘ/i(2΁҆�2(�i^�e��5�j�c���2R����qpd������"��S�8,�27'0lH��|�,�F�w9��{�3�w�������������w�A�p{� 	$���=7���V�7w`|| +���{�nffrI��7wbff`7�݀�� U@�U@jT�$> �� $� 	$�I 쑶	{;-�W��UoG�����!���s�Zض�$ԝ&P��ed�sG��ʤ�U7T6Y$�Z2�v�+HW�sު�]�c�J�Y����w[m�a�;��_fer^I�w
)|� ���3���W�+8��k�'T�E�j�u���J'�UuБr����6���Ν�c�`쓭e�ֽ������%T5U]���G*��֯dQ���d���:�ͫ��uG��U�$��Z9ٍ�M�/+3��=���j�m��{ټ!P$����F�)��V[!��r+y�̮{۹6��d�UP/x1�_&Ϸyi�Bm�sj�e���Qy®�Y�n]�@�l ��}K�]�I I  �H $�����rZ���-�ZKn�3e�_ �lv�%��S*��K��;jX;&�x�_+;�ʹ�r�}�˻_�e�T�d2����k���U7T$�I8�ef��V���UT�V,�B�[W���m�M�~��r\�]�̢Kv�/ܾR��2��z�_!��̮�s:AN�&�do3I�9�]2�7�> ��Q^�q6�|�lzA����)����칚�km(3.�Y)���&�r���(.��3,�[6����_�V])TP*���tRփ(���i��	t�����IS�������f�v`w���uw\�,�ܣ;�3'L����ըz��mRr7�T��rzU���X��K��yN�0�_�
�G%���'�U�Ǭ�Ϡa��,[���Ѫ�kvꪫ]��U.i�l�I����VK����f�wf`�#�|{���q� ��f`0{�.��S��^��)���&_W�N����)9���Ax�t^��RVػm�A�f�9F�Z�O=:��K�v����4�%�d���5�=�}��Ϭ�,���͵����eZ{~Z��������=���Z���o�]��|�%^X#�L��윘�lX�ɁULC0v3 �s�>���L��7rc�Ov�(����8��Lݙ(op5�ך�\�:C��*E,κ�Ԓo2N�˘�ܙ���^���L 1l�� a��O��ћW4���67�����2�$�3��O����ԃ�3�dco���}UA��@��\��*D�b���xXtNo��}.�Es:�9㪪��H�P�x`k&�'
@��c:�����Srg\�=�z����= �J��P�����i$G�z���^�����$��q��_��b����V��o1��9(U9s8����Gd���lZJ��uɲ�\�G�Ǳ�fz���\\-�)��Lݦ]����k�w�*���AB�0<���1�����z�3W�MڄZ�8�e�f .%�|��O޽���2>�7dl�}���v�ٵ��ݓ"�76������i���}R������9d�[�#�˭���+ެ�\�����n��v]������`Q�gl�ŗ�F��$��oF����u0͟V��<0׋����SL�����<��d;�/h9���k�h?���S�T�F��b�O�ƫ��Xϱ[����K����8ޞ�̗�~�j�jE�Drˊԑ�Sj��=sI��^�*�*%���G�8�Ǣ���/��e6↪����4���|T�v�s/	R=r�&�c��S�0_ݖ�k��˻8�w�^U�M�|��4�#���=_��mxd��keGW�	���ݣ,]$৹�_ad�f����|0�ޅ���	���̚I�UK��Ù�����r���5s�*�ڭ�*���v�d�h��U� �F�7T�mu���｟��������̙5l�������ٯ$�G�ߟ��@f3p ��������Y��S�^�z%�β�jv�f:�;_w}�I
�!d���K�t��np]9ga7c�3 �y9�$����W�{�[�R1M�B��HlU@�~ٝS��f<��H�o0`Y�=���a-O�	��2i�����=r�I?xʑ8�'}4��b����K��ы��S��o67��b=7/s0���~r�������T�^?=�����n��EUC7��B����(S#� ܐ���b�,��H��W����G�wH��?��5N�)�Λ�;���Xvyv�o(>'_0�����ٕ}�M���V6����i4sr��t��jkd�f�����}7
J6Z��C���s[t6^w�����s�E�}6K3{�:^ifk�������0	����GO>ff5�X�s�i�S��H�)��`�ǂ�.E1{^�ﻹ�^�t���߄<��������E��M��0�,{.��	 {T-U�cЪ��4\�⾘S>�\��1E�Y�0�}�Z�|aI;�~&:��}z��UԠ�r��nǁ����M+����Ov�f7H瓇Z^)&D��-�NGDI{	�RS3 ٞ�H��W�r�2:�����6w���¶��*��n�ܩ��lQuÃ���[b�g9���Jb=QV�.p�oT'N�T^����(�p�e�_�a
�NGu��ei��s\�߂�z؅��C @�v���mݙ3^�ė�����Nf���ג-كu�2mF܅��͹ۙB�\�$�7uH7]ȷV�ٽ�߇� A	��teENR8��i#F��EO\M���{���d�m�k���x_���G�wH�ಚr<�3K��z��C��r�O��0io)� ��.6L�G��Cwh��{DioT���%l��E1x���]s�����\:�S��M!�H���� ���G�;CK/��VM�PB�d��
��+B���X+3��z��g���$���,v���?'UG��B�:��w�ݽ�����x����3��MڄZ�8����y���z#ˉ�+`�.[М��|��כD��>*F%OPaE{B�5�x�ٙ��f��`d6�.����$a�ۓI[�6چ�6�˕r�"*�On���0d�T+5���v��&�q.;2�\�B\[�����5�Z�s�wI�"q�w}$�=��Ã6�f�S����~�w�7M��J�cT_��:�ę}�xt��y/��s�j6a�h�3��$c�R"֞�û���PW��3���I���q�s�Q�y^ɾ�jH�7��ա��P�
)�(sG�)��#�b���ǭ�VţBY�w�[� N�5�~<��n33h37�FgC�<�7Jz��n>�LU��,�!W�n�"~�ww[z��R~"J`f��:`*i)~.����f�p���,���#,z!�����*{j��=Z٘�u���JN�W�)A�>�"D"V�yY�\ֽ�֜m�z��(�g��7OEn�_����]��b��7]�;P+*��x�5I�M�}w��5t�pT%�CTۦi6���Hl"Su�l�������������xx��v�����z0�E*^��
��5\U�V���*�NL����TG�6(�8�a�`��H��n,�(��eUmc4/0s��͏��I�߸ȩ�/O*&��JwÉ��;�fX�Z��kڞ���ޅu;qǻh*)���D
��q��g`��r���/{fU��T�k��N31�)"�ID��D�{WC��^�>X��V��o2�w`f�z��f�*e�=�E��V�9��Jr6�7�����KӍg�z?֑���zó���O咎^UPPa��ķb!P�S�F�i}"��
�S��~(w]���u�P�Zws.E�{���D�9�{�1�u�l��`[]*��JH�N�o(jI;M*ӥQQ���E���m�l�M'DRc��L�Ȳ�I]|O�n8�d�:C�Գ���S>���+<P�7"��Iۥ�/]��dx�
�`������W����j�fO-ēɦAI���m�v>�J�wݬ�D�?�&���[�Zl��H�)����~��w-���'� �#�9� {��h�bY�P���q��Y�R1~~��n�`�A���Q�2��C�0h[��)��}�T,�7M��<i�����>%ڙ/�@ͥ��<�d
����W�&sr�����4��\s]N }����RE�)D�ĉ�SȤ'j��f%���p�o�0IC����P�ԶM%x~ 5&L{z����L����-��$�q�u��E��p�]t�G0M̥7NBM�V'o]�s��I�M��7T�t^�����}�j�)J#�I�ޱ]N���S�0�7��������8�,z\`��D�d.TС���D���z���"hog1I�ұdN9�@�OQ�"�䖀C9��ȇ�[����� �c��w�����N}�[���^߼S��{�ʺ���jt02?0�=����Lq���2eU�h�P�!q�`6�|2����c]�հ�ͫ{���χV~�c<�EC�[���_W��8��{���lt=��, QX��j�ˮ�t�;Yv��hO�eP�s��M#�5�^�Ϥ����ت��H�)�Lɯ��G\��\zU��G�#�����6�&�fll�u�Co��L��Yݨ4�b�L`���`q�	BP�5�|�$��0��(*���1��3�e,X���VXʔ`�� ��b#g ��z�:�<<�����/�q�kLØ��S333333>�̝��љ��f 	$� ����s30=�A�bI!;�  �$ 	$�>�d����{$�H�݀��6rJ۹�I=&d�����H'�L ;� e�� 	ws�R�s30�H I	���$�(r��Z3'j��-L��v�~��ɰ���[y�.�;��ؗT�K4����^�Q}��H���&���]Q�e;��0�Ks;����vD���=�T�ѲI&{6�u���|�'6�G��]�X]���"���w{������Ԩ�h���r�Q�e��n��7x���9����*��$��9ۭ���(��V.��N��Ӯ�1!v�v=��\̦��7.��U�eݻ$��s�F�i,��R4�.��ʶ΢wv�e�@�ْ7N�'��6���{�7s��U��ns�w{:F�I���$�O�������+�g9�lgm��˜��k\����:ړ\�|}u�w�����n� �݀�� nԩ\��H 2I �@�����_5�6�.��`�l�m�b�a�m���WkM���.\��D�8l��WK6�\����[��[uRRؙ�ȹ�*�q�߾����>�A��Z���j=�;R�(a��̽$��z��ުD��!5F�B�j�;�)���R[�ܔD���$�n��,�ڦ:9#UJ�9Г;0�n�O��]�w��)�/�R��3:(!����pB�16�p��(�x��>*���D�aN{�&u�;6t�ff a�o���g�M�2�7&��bI��;����5��^�YKv�V�a�6mSۖ޹���r�wd3�-]f�V v������}��~���.��7f��X�D����|�����W��~�ۻ��>�T���D���|� ��c#�+4����~8��z�=s:j��[ڤD+=Y�YE��N�0�W�=a�M����l��Ģ;��MM��z?uߔ�US�e'Չ���H�-�	}�N��n���/9v����~v��l�D�ʉ�g����S�3 �z�c��TR �D�.������ڦ.��ffv��uL�2�ffp����%$�x�v!���o�o���_�h���������}$� f�|a�f=��QN��&8���E�G�[�fbǂ_�X��^]=w���q&K�Q�ۘ�/��f���<�F��hdYW`����o&�z�����/߹��y߾�[�߇6����2:)�,��h��w&{r�&u��� ��>�4+��B{�; �T��﫦;�	�UC�U$ȝw�h'�mآ���ʣ;��'l���?M(���G9�TYvNϚ*�[ N���޲�(��0u*�̲/�O��IS'����_J�"���3"���Gz�
_�&����7�o�u;I.��W�Fʗ�FM%p��`3A>⤛ۗޅ��Kl�~��"�.-�z��M?��z�^��fcҲ/RDqm�Z������Ui�y���ow��l�������͚o33q4_(���R���2�gC���B��a�Y��A��]�B���NO���578Õ1��͉�u䐙�w�M�ij䙚lITuj���x�[u%p�*��k��9=�{�y���*\V[���B<���xt�8|2C-���>�w�:ɳS���"�)�S^��i���e�����;�������f��ڭ;�g�+�v�333E�$a�D(����u����V5�G��q'(���ez�0�T�gx��UUo���G� I��f�K���:�2/-oV��ܼ:�ԛ66�E�~��x�/�<���=�2�bVFy�����:��=jH��Q,6�=�35.<��ZM�;ɲ������^��v/׽}�s�>�;�\�]ZV�5M%p��9�dw�W�3��[k���Nw������%��O��ŏ�>�1�Qx	)��>�ow�f}4��UW���x7wd�wqI��wӺU�k����T�C�����$���[�&wZ�7u�{����qQ.�	#���S"a���)���IP{�8C����#+�컻�udF}*˒�F�=M%ƌ�dڬ����uLߋ6�� u�v=���l=�E5<|4��|�\�,�/������Rr<�>��7VX�m��2)�}�]*��YԠ4,�{��nS�=ü4)#�sМ��}"}d�j�2��f�{��3�-S�;�KqԡDD�+Ŏ4aB}�~#7I���o|>���'��\��[��oU"͊;����A��� ���}3�o��~������ͻ�K���La�V}�X31�#��y�Hȥ(��8��5 ^�dq�\� x��<����Vﻇy�i�4��w�Nz՛u�p�����:�Z��ٌ"u�'v�ޮsrξ�l󤽝�p��o:9:%�����TY7�ռ��lxQW�|[�-�3]\��A����Ω��uD.�l{Ya��{�3�����ed����"��x}���-f!0�V�'�?]�uoY��	�<%�[����9y�QL�9���U-�ܟZ9���႗��=Jo���RR �Deǽ��ޝ�îǱU_�2� ����̽�������i�=�}S��þ��'#OA/��&���/x���/s#�B�YT-�,�٪p��dS���x����˻�|�	Č���	7'c\�=����^�2��W�#
�R�d��L��عV�Y3�"p���ә��}�M���Y%w���K!2{�r�&8q]�(Y��L�]�������=�c�۝i�&�Q4i�R%���z/d��k$�v4�?��Z/��jǁ'��2�����C�V[b>���7�ì�F�Iۺ��J
�"�3�E
���dZ0�_���{.��������"�ID�Ď�j�)����^�Q.lq�cռ�I�3n|U�*m���̫J��?�����j��M���/l
�����������{��i��ǽOSI"8��x��:�mx�x/jq�OMNo=�C�
�n�3�O
{�e�#���#K�)w��.�� ����7�}ٙ�Xtǰ�i�=�E3�gM���=�vr�z��G�<@��}F����C��Mݨ�~�޺DQj�C��(� ��։w�=9�i6�˻V�o^�wvM5ʥ�)j%�&b7�����j�a���k�M�4F�9�&�������$�ܕ��Z+{$5��^��P�G��\Q���6
��-01�����c���R��`7�I	3�h`;J��37L��h�����>v�˅�>Ѫ꼂�uL�o=m�:J^�]ש�(�Rt����?F��UB�rX`6:(� �-�D��``n��������^i�l��wn���1�P0Nz���<�rC{���P�}hʤ���u-J[&��3�"ҭu���(��z�44	���쯾�s���6��Aq�>�}r��[YB�+��$~��ԩ$F�2-\��p)����w�|��P�������9IʏzW��_�gP+�����y���`�w�$��iv��-�Gv�n�6H.�ٹA����r�ʙ�!.��jI�M�R�rn��7����%�[�Ѱty`�utؐ0,�lU��o.j{������j�|̔v0�ua��`��p��}��ݫ����#�y�I|  o5�}�1ٙ��-l�n�gE:�Qb���-�C��JL�̼���707F��^}i(�NҸ�N������ȭ����Q���9�b����aO0#��.�w{Qo����f�V�����7M���y�(c
 ��qmnr�_���	&��o�`��G0�دU�w�F�e�g��MP0M�LS=��xP���g���b1�]��?^k�q���4N%p��]��3 T��S3!K��矠����$ir��[�p���\��;ok��ᵹ��w!�����n͕���uw�\��9���N�͔�I���ίou���s�� 
�������;���dZ��)a���6#KzU2l��H�j(���[�Vw�n�T|?=�h�kz��Ovdf��"8�������e$��xW���"ȁ����U]��k]�ژf���{��=��~���lٳS؉����^�o��/�����<�Wwj/����n��*� �.,����y���|�^�m���b����`D����%�M���*A�O��Vƕ��[���[���u_�@���0�wϪ��zu�x��\�GR�IS�f5��h�~�/��HH�����Dޯ��w���w��_��hwfQ��ٗ��X�uf�n�W �<B�FI�f+DVF�v�'߷Ͼ��x���/�2��[�U&��SLL�)��݊v�v��@��׋�c~�d�F�wNU�tD��H�L}�Ȼ�0M���(׈�r��&m,  �l� 7���ul�����w�z�j)\����i(rǵ�3S̛��&����׫��Lw�:�ت~$~������ED\$���U�>���B���bȐ�o��''�̻��QS�y8�<��|����&�u�v�O��!��D�:��SN�e��lS'.�ݭ��9����H劉�{]%;����^���u軺�[30ݎ��}�b�M"(�(�ҽS=9�[�����BeV; ����`�� i(�}V�{��נ	��|Y�����7K�9"���m�I`�Ն�}$�,2�	��:�'�t!F�@�@p$8�������%�����gB`>z��r��M|�Ɛ�DԧnbtX!c��h@�pv�"��o{���̛������wv{�l�� �d�� �� �@��I��������� 
�e/��d��{3$�O�����z����? 7w` ���f` ]݁��o9�$��@�H Iowdm����ɖB�l���')�r��ւ�KU��9�N'���T"����g�o��n��g�ϲ�v�﫽���N鉺�Ȳ,)uD�Q$�{���$�6۾��{+b��Dm4����E��Wa��oO�l[�nb�����mt���j��NɻVi!9-�ή���l<����7�f�^ྨ�[������y����qܫ��j���N�j�'m�����.��ea����I<N'��F��ɫk�k��I�uwm�����a;��1-WMS�I�F���J���ߪ�oM�d�J,�:$�W��]M�{7��h�ڱ��ݸ�+����>�z�tt w�@ �݃�W��$��@�H I �9ޫ�����
��e%sH���ٻc�7[��-�ږ����\�inK5�`�M�����s��Vh果O[8��2�{�`u.�9��>˕ۻ���n�������Y��i^��Ԓ䒾��{+b��H�F�g[vk�ڹ��MW
ӷ.K��=��!��d��;�;[�Z_|��d?����T 0�	����D`�& ������@�aS �;���v��F�Շ�+/yI��t�m�����N�s�7H�ѽ��o�cs1�ͨ�D�<��;{��ˡ��ޞ�_N8Q0�T]ɻri�ޜ:F:H��	�N\��^w�M>����S Sy��'�W̳�#
�Qq�S�/O*�RЁ'G��2������t��7��WU3��;<�W�������3�(-�D�������3&��ܞ�I�UjH��(��� w�fϋ#Hw�W���&�z���(|����jZ��30��[�lN�k��ᗕH�S����&��òg���s��x�m];q��^���v`a��{ؖ���I%J�-������O�f�0D�(���tq������.��Z�<�2��PQ�kޡ졇�8��T����ݛ}����<�?�={HƳ"�=2�=e7[�����=UGt���+U���$�i]=��oL�gvlM's*��g�ng"v�;�!;���ӳo$[��]����er|{F#[_�P��L�-�]���a���0��e���u�/�jb#���]��4���b���>
||��f�����ը4��yU���O������Y���ϫ%j҇q�I|0�{�������ø�]�d]g٩���J��������k��,̗�KE<�de*�.�{;��q�ޞ��*R6������UT�'���!j�3�1.����ʷ&RNz8�������`��Na�ʩ�G�e�����0�
a� |WD���x�)�ﲻ�컫��QQ�'^���#9YQ[���b���|p� ���)6�_Ia�ܚJ�Q�r_��˺{���^m'����e�n����t�G�a)s&�ڿ?z��%��m��o�د>�(wD�d	��Pc3e�t��R)�d�qE���~�iYU�.Ja�9yȁ�r�qe�g�o�32斛ZA�Y�%��gIf�,McU�|���N���ӏ�v��UA���2��G�/�Ë9�i��uQf&�:,�ċ�d?�<vA��Z���x�+-��<�F�NY�e�Ϲ�"D".'�j����8�Gb�0�9�2
B�t������Uz��I�F����nΤa�6EOAG����T-��1��c�Yhx��D���Z��6\���߾��wr5$}��&G8�_�J`r��$�)��ﮀ���F{�s-��$�L�#ܣ�.��I7��]��]&e���tA�<5�3�z�ھ>-+s/�߽�\�>���-�B�DnSH��^��՗�d�b�/�?v_k��c&�I�ټ���OB���D���g*�BA"�TS�x=a�	+,1g�����U�z��&v_zG�r��\�9Ƣ�Y�H�-�EL�'@���W��n���/9q;^��Z)��STQ�s��r��ҝ���F%"�F�x�ÑvA�J� �{��T�̶�xx�)��.̒閨 M#������oe�q�V�A�=eժ(k�,�ط���F?��S�n�c�\9�����-ɨa�<���+I&c> �%۷�,s�:�9���Y��]������G��VxPn�k8����xs�r�F���Hp��&�;
 �Djڪ�g�����U�y��VwU��^�ӝP��D�"�ҼNJ������7uܨ�ӡD*['=��L�)0�t�rN��SsrT��ſ|9�;��6��\Fv�H��r��*�K;�
�(,MO���ͷ�CüG��L%Ěfv_�a���NV����=u^���Ȫ��	��� q�"_���r�̻����]N�K��A���	����.ه*���ʣ�I�ܾ�(w�2��%?��6
�h�{�}{I׋$�V^�N33=K+�YnR*d��1�<<�X���oj3}��ws�w�����r(ʝ�C��#%0]�K������ސ��4D{�M���[3X� ��Z���k2[�L��&%Qm.Q�%���4��xrь���)�f�i�;R��1x��ժ-�m��K&���E�9�ԁ����j���G�����I��1�"ŲA�)���a����P�t͙7�8�I�M�]&9"ū2�-��Ͼ�N�:��۞��A��; �<���Aow:�*���}i�;C��a'2/Ae|�����u�UU{���)��`������X��{"
+5�Ԋ���Y�ٗ�R6�
/Z
�PX������^K�y�|"Ĭ��ףu1#����I�R%7p��}ҥ�U15-0�#K� q�"_>$�ʷ"RN|mR�H"�����~�I{*f�b�&��J���������%bbZ��/ʌK�+a��� ��߯=P2N�Y�5SGQ95hf��v�?�wF+���˻�^:#d֩,��r�YU�.Jvs+�	�#�8o.��f�n�p�٦�I�����N�rR�Q��μ[9^�uQ�f��j��޹��L�$��K���t� S�pOT��]-x��:�&���A�t��J)�΋��yL�ōXY��H�1 �GJ-��E��h�_l^�ET������5�mWzK*���'E�8�z��e�{ݲ�Ji�d��H�G�9��IAp!�^Vk��2�����9�Uk��q�D�d�ȾY�'=�*E�t��tELD���w�;35����׾}T4�]��d3�Gn��1��r����/�C��,�R��uLQ�x}]�4Y��l�M�z8���M?�a>��Dc��q���)'2�"(�vك�a�������UUXy�G�G1���I�X�h�s��������3�~��{q���2��lҪ���;b��-���1мk�e��{�1lwx{1eW���MҦ�1�����0"�@3�f��������{���1��æN�<  ޼ݩ�n��-�� iY>�N�qD@����f �v��/d���EzL�����!�R`�8���71��6���31кu~g��>r�YU�.JE&�\���&������}D^@�����_��,�Y�DV�o.��4�7�}<9h�P��)ܓ{�T<޼t:��/���$��GE8�z��G���G=ԗ3}���`�A���!yT��3�Pka�#1>Z���x��(�����d��9�d��q��eՖ��xs�r�Fd�&n��k�����q��pC�IdSA*ݽ��P� W�ux��-XA&��}x@���������nze�՛[iK�7v�&�hw�L�e�!ՠ�:Gk����5�د!����h�W0>�Og��N+�FU�}�I�-}h#��? ��@��{��=���y�K�fb�$r��M�o�@��30_��#�ܫyQ.dxҏ9v�J\3�_�qFi�A,��P���WiMCP� H�W4P���U�1�6�v���w�V���uer/S�UAŹH���R����pH�)�~�E[�@�|�Q6|+�y�}#��P(��Rh��4r�q5��ytz��ٙ�y���i$5���4�GQ^�L~�����T�P�
V��0sQH�RA�:˫T_9�u�Id����t�j9;��30x��T\�H�TA#��K3��Y�/wsu�z�x5����M�Z���?>g��;�Z�8��
��5}�J�L��n�Ę�ݻ�6�w�·�n��>���0fj���-C%��;�=�G�Ԓo3����$��w��w}^��wl�9g�2:΂��� �$�O��i��S7�2�4��w�����&fff�`�xf�������Ff�UB�r�^X�����	<v���ɂ;��1͓ۻ���:�����fc�*�~����8n�cޗ�T��~I9�4�0��m��N��	��c���n}��t�(+}<lZ�$���7|l�i�fa� N�%���8���۴qj'ޤ��#�!"�[߽��H!{�c��ر=���v��Z2�d��8��r�Mɱ�;��a\���d��^ �����r�� ��|�ʅUZ�eސ�dEe3Q�m�I�j�xr��`w�e���[7��CL2��Wy���HJ��cm��Ѿ&i4c�o�����$� ٷ:QL�5�6�L�1I]�М��ۤf	b�S�|��"p�b�""&8��; HI� -��� �"3��� �wwwY���bff`	$�|������nl��$��� I$ I $��=�y�ɲI3wv �H�IUP77vbM۸��$�32}$���e�f 	R���� {� �I��9�O��߿~�\����r��T��]7$�����{���wUN�nw���R��|r����7�)fgP�Ȓ�휂�ͥ7E����jܼ�rI$��Ȼ�^�n�]���tI����=�T�%��I��8��
��2��N��&�¢�ݲ"��&�����-e]�����f�ٚ�U���ޟs���Mo9���f�pnq��W�����d��L����t����+�q�}�U����w۰.�7y���U+g��jveTjpC*�e܍ѣ��a��N��a0&
K{�fg\�}$i$ٜ�t�R_�?�?g3;l�ˣ��la6v�ˮ6s��hj���,��~�߀�3w@�� �� $ݩW�;�  �d�I!�������k�mWfY�d��"GJ���5��cU�k�`,�ڐ�is.�Z*S�l�[湻!G�)(�%��cj��\х��kT����.[Wq'���������5����<��ʾ;UET�7�)fgP�Ȓ�휂�ͥ7~��߻���bgx��!UA��.�׺Y'2�ʵ}�&���ɻ���ii�#���%��u�
����:9(�ɛU*�m߻�<�  `����2��<�^���-o��ߞ������f���O{�6쫼:sa���W.{�]�7���ȳ�;��rɺ�vKv�mf�L�2_\���g���v{�����b��TC�����P��ᗊ�F��}�0�rnS�-ک�h�c��q��sԬ�G��k ��*�+��{3h�mxc�M���8�!FɅ�O��������)��f�I��>q�Rm�-����F`![0�N��ڢ����O�>��H�s�o4�z��5?GB.�I/�:�+ ��\H��6h�\�$�jN�gz�nf]���A�7)� {�4��3�2�{��U�u�Hx1��ܩ��DB��D�:NrH/gG�w¼���#;M����mS'y<Qp��ܘn�V�&����"AyH{�>f����;ʢ����$��_��f�����B�Mם�s�m�j���a�jV��y�@�:�b���$�%�}g�W}�^m7y-h��k+	���g�>�{��w�'���0�0!����*�����̣�%�����)�M$��^��)�#��&"�z���V<<'"��14bװa�VfM�+����?�ݘ{�����9p�S!���6��A`�g��Ǉ13S��[��K���F�x������Ū-��Wy��M1dYÈmWۜ��C����
j#I0�(F�0Di��lͮ��yԳ;}�J�1GIE��2*�����3��wp��4��$�$�O�� �]�ܚ$�֒M��x��k�m��qH�9T{J�(,MO��2����zt�zİ�ƛ�}xm$��i@�H�C����Pz__�G�s!�Hf�)ŸA��r%$�V?��цk���n�;ޛ�xN�k2�Ն�i�7�;��vF�:�Hv�x��v�X�%�f��-1M�4F�9��̙�29�,~����x�D3Gt菾���x�f��{G?�%�3�qbm���D�6O!�Eb�34��z�.]����*��/y�'\Q'"����=ll$�TY�ܴT�D@�ը*�o{�c9ᙛ7#bw|E��V��zj�Œy��9eT	xcA{7�z��"w�)\R�wDVx�̂�r�\��Ox�Y�36�$�5�xr�V�1�;��������2����';.F0;!W��c�*�u7睗��8��D:ANpxt!HQ�)G'�AV��S{����$ISڍh4�[3����9��dP��|Wܺ�TMF	4h��'ƌĘ��{�D���I�R-������vt�oy��y��݄��+��y"ݘ0v�}�1A������]�N�t*����A��wT�u׽�#�v�54mnV���㍟!y)�?T�7	
�e���;fZM���ׂb�4�ʫ��z�t��1��cHw�Xm�%��L)����6�����}�j�S�Z��k��CZ�x4sȑ�G��$���oA�tZ�z?G�6�ʉ?W+Խ����#�!��Z��UT�A�Ev����"&�AT;o����5��y��vwg�����$�>�'k��rʨqr]����!����#��Iۢ	tF���Wkь0;����`�G?��e��X���X9h�l�A�=d��Z�F���ꘈ�a7��%�NBi�"�$^�c���X�AƆ��3�*�*�Y��$���w�q+uy���_��N�}76"�z�4`��s2���7��Z��v�ɫ��sj��W�q��t�ʍ���f\���33���{(���f *��7y�<� �p3N�t������[#�kl�X��	���^s�C�D�W� �]�T#�>���r�3�Q�>�ߋ��$-�"}�����Pe'e�Ùns0ș�
<]Ď���fa1��7�ޏL>��u�^�0�ĳ�N;K���L9Z��NN��d:%!���BuTG[Ԅ.{�1��tD/uNtt,����Q��rc�@��pUfJ�`�sg=�Y�v]�r�m�2y:Uy��*� �ܤT����С�ܭ"7qAT;{Y���g.�˝�ڤ�J'1<Z�~�iYU���Rh��xZ9v9��h���v�7*!8�d����9�����hݝ��s������ͣ��YW�:�kiӦ�t���f��K�*��Ti�e��	QM$�-*"K/����v�������Hs|>�)�[����ï��`���|[DF]� �4��͟u{|��xrb�w/�ˇ-� ��)ܒDu�V��9��o��1�]�.C��5��y33 ap�E�Q��H0����5���ͽ�-�����V��s�����̫����1�\\P��	�@�Hf�M��=�j���`�u��\��*�Ü�`$�<���7m.��1ҵ���9�p���{r���mA��3k#}�~��������s
v������ �NE'�33�<a�_N^6��uTG^BС����4�'�I9���ڮM�Z*l�$��pU6��6
�h�xe����;��"���ǩ$r�ݽ՘޺�L�E��Xu��"�]���O��i�;��ke���z~�'rZ�"��ӷ_C��A"u9e�}�ƺ��VVT��D�j3S�UAŹH��:����Wm�V����qѿ�PkO�(���`��A'Gk��x=8(�d�Rh��x^��NWq{خ.��fe���9�ir��E�X��~<9�S}�Vgv]�G_��0�f�2�Q�s�uޒɧ?4��.Zތ#�H��H� �ܤ(���w�+I&cƏN_���e7v��`�A�aG23kv�}O��ü4W�=��I�� �1�}$�Bk�[�fǻ|v�n
�5�ͥg
L�fJEU��k�U������f*E%��Up�~�ë�u���2����]��o�V�ow�I9�z]f�5n�Hz��šx�fR�zMĎt׃w�Ogq$�����f�"�ͳ��{W`�}_|>3^)λU�����<��ND�i ��i�{�ޭ�u��$��<A���6k�!���-0K��y� ��|�(w��lm�3������׌ُQ��>fc;|�O��fgixҸr-�EN��"&�AT ��W1~��ۻ�����E�t���Q�^��*�Q��SW��ϰ�ل����/�E���0h�`��r���K����C�� OE���Y^�
fM#��R"{U_���f�Ը��J��R^9�m���dӐ�zK�Ïs�����i�$} �nS",�)
� ��xyx�QU��t��T^�k9��lI#F`���w~�Y��= �7M�4��T�ݩl�<��w5q8�os�,��u[9�Nڧ�-�s;x�����rv����a������1fϬ˪��q\\&2��ff�$�3*y��
ͺ��}ݙy�#k`�1�*�At��t.�s�g���e�{�K��D^f�l���m rS},��x����Lʅ���'1���
8�Lr�Ȕ��S�� �Y9�;޿vz�]@�ʝ��j��Z��\9��GI�I+���^U�4�:
�,fR�7�L��&�r/��*����Iw{0�dh5;GQ9L�ԭAT;{�3���ðc�!\^��]���荓Z���6�9ET
8�)&����k'�uĪ�G�����$x�)��v����L�4��ABiH��kr}BDP��3!g&����03�;z���۹�%y�s%̻��y���̤��e���W�׎�{���r��UO��gNC���[(�Ie&�l�MR��t�sN�d��Id��/�6mTW���f^�q�0�k9�_<��:˕É��ٴ�}ױC�s%X�A�9�5�LH�}(���Z��n셹�^����Z��t�Z
��VY7F��UDH5�t�Um7���
��mʿk�����!t6nv�g���v� ��.AW���иs-��D��e߭z��"�%���G	�6��G*�cAI�������'�VN'Y�ۑ)'21�<Y|������?Ӽ}UUU�4IH�D�2MrHX�
��=��0����|���+>#�<�˺��DE�r���<[�|͙G��W�ꘔ�N�0������r	�PUۯl�A�o��� � �#��P�����/���@2�M*��D(�	�ءA�"�wv � �"B�4��,)*����(�""�2L� �UUA���$�'� E IPP@����$A�D�� �FQ&P� `eA���B`��RH  d&`�DT	RQ�@��P)�@% D�RR VU � ��a!F Q�!YHP��dA�$��H���(A�Q�D����`�l!@��RIP�� ��T�&U��`� T�AUYD	@RY XQ�U$Vd�b � d�R �Qu�"��X�� !Q!H0qTH@%&O�~k��p�{���*��(� y}}7�����߇���>���:��?����r���Z����� ��G�����z �#�~I��Q�X����`��`�`���������A@?������w�6����:?#����������/�?A�� J���J���! �� @� ��0����3	B L����A D�AJB��
H,! ���H!"B��$	,,!HJ���B L�AKC �!+@�,!	P�2� C R�!, HB��$!(H# !)(��$H��J H���������" @�$�,�H@���K
��J��(� 	J����@�# J0�*BH�
 DL A((BB+""���
���  '�B�������
�B�2�
�, 2
0 ¢��P�T�!T�d�R YUEC_��I��1��� ��������M_����p}>�������}7�� ���o_���ϧ������߻>����ӿٟ��/>��� ���������|��_�(� �A@9����0���i���D(� ��X�3�F�/�3�����E�;Ѯ( ��������A@?A��?�����w���S������?�}�r��g����s���� ����������}_KX~��?W/�ϡ�?��=�΋�����y��O����^�D��?:;��ڎ��*��������07��9�����
?OO���������(+$�k8sa� O#��
 �� ���)�þ5B�@b�ۧ,gP!(viz݀�]��@R��+4J��ѭ= ����t��j  �    �%��Q+[B�!A�Xi�LM$�-2l���ѦڃF�a*�kh[6��ִ��mh�ƥ�  � )R�����}`W]�3Tc`W�u@�X."����=YH5{:AE�Pp�[m
c���,ҕWm�\�B�s�������vsSm��[+��滮��rD��t;��^<����y��r��M�7�R.Z�x[���z=���U���[^M�8mu���:�ƺ�[N�xS������t������j]�nr
�(����Z�z�����nr�
A��kt,�P@��k�5����8�*-jp%�k��Ӡ�������Z��'
ڠ	� U�;:P��A�5AY@����:��T��p*��9����G;p4Cvup4��*�a,�fV��4
�Y�G �C�g@R�	 �:t���:�(q :�wp�P	mV�
��4���Nt;��3i� �Ѫ�+h��
�5GGT�4SV �s���@ 
�����tl�3X
�5�5�ؓ+@�����Aq�'5�     �J��ъ�J��hh	T�4h���di�1F
��R�Ԓ�  ��SЩQT @ ���II�=A�A���T���Q�  ��l�2�?����������o�Y���h�Ǚ��%(t��r���PX��J�^$�j� ��P����G����o9dU�*���qIc�mK����qn4m[|��%/��L��F#t��bR��;�8���\��E!f����ɏg�����)�+�s+��Q%�ϙH&HL��[Jh�8:]bz�^'k.qg��v�!'Ę�7H�6�LO�S���ꔔ���Z�N�Yj(ܔ%b�b�b���O��R�2T0]�G��e�.;L��Ü;3���g�K>)�-)�Ϙd�|�n�Ic���%�%�K�؋)�)�:m��mh��Ԥ�
b�-�R�mvڛ[�RI4^4����&�h�;���JJd��iK�S͜����ϽȬ�	e���&#m)�6�Y�iKGx�M��e�h�%H�,�4�d�TقYm>(���ÌJ�O��Ԓ�4��lnH��-G5��+Q,nZZ"W)��ѭ����2[Cjc0�Zh�1F�`�l�]c�B8q���g�ok�SblM��6'�&�؜��SdlM��W��Yzt��;Ȧ%(�sD�O�ba)���k7\պ�K��>�%*���"ė������Hr>=�S�G�'^�=�E�z3}��Q�r��P��F9v�ɚ|�1λs�^�of��;ɵ6���R�	�X�q�rn_v�L�O�����EE�i�i�6\q�����Ó�A	���+笟_a�Y�/rɍ[ۻE��}�颢�6����|B����s31:ͪgQm#hT������z�\�Xr�6���ƛjz�S�p�Nmc�}�f{�2�7�i����6M�c�F.Ӭߗ-��Aw�/�%���4�b�M��T}H�����d����e�}yb��^P�멐�'���S�Է- �B��y�*�Eb���w��B%��@»������B��zJw��|�n���K���D'-�>���cӲv}]���z�����u ��^�z��H�/��u�W��zu�Ӌ�T�ˏy�xw�{�B4�y	��7N������G�_fZ���{۾�_+�}ma�K��|��#MgO����6)�Q�@����>)|	2̓��1?��}�J��gT��l�y���y8�7�����7����^�xTk�#�:S"J�$���z�E���T��zE�oQu�����>������ub��x�#�C�����Ǵ����z���o=����IǱ�B�9����I|<{�������=�?���l���M&��G#�P�N'�L�f�w�V��S
��ﺟ4Ek>��}_}F3+�;�:'�L�꿭F
����~������I|�=a�!w�(ZY����Y����_Sw�K�6�>��WaE������iK��6�S���N��$}�<K��k��K�l&}��|Jܔ輛����Ǘ�=��2K�����
D "�F*�;4�x��)���
���5:���j7B�kJ�&�
��i�}���=��������y����5�N����:7�z'
Qx��D�a�D�@���/L�����8,pn%x:h^ݓ�+ݺ@)�^����M��x��~�*�H�w�����y藌[{�=����Qhй|Y�l����R�i��[gjV�Q&��K)�5E���ı�%,EL��Hi�8�fqٜ��q�鄉�E�ő��i��)fSL(�hj4��AHP1�[n�C��OK�\cffg'�q��+=!H��ٞ��]�K|پ��u���2����.1L)%%r[m8�KR�D�K|��RK8�+n-��#�㜜#�W��,,*Q�|��(bEI�m�.�|���Z�b1()RC�E�i�aN)�ϥ����>c�Sd�$�gb��j>d�-�:ԥ�Z�r���-�-�%��Sm>[jc���
�$&T�e6F�l��:��*HO8��)l)�ێ0�N�֍���(Ԭ�*V�,�%�����b���cF⎛m�|��J5E�."�L�R,�鏜S���\��[O�bUm�_�FIARE%)d�4|ԑ1qN#���-cJ�Ϙ��;f]g�+��ى��0�R�b"�pIK��d��&J,�.P����x��aŗ3��Y���6ю��C�Q')��l�I�ioN>=>��#i6S`�����ҋ6��""dH���"N������Ne�\�ՇN�7+ARąJ�4|�Jb�6�.H�j\��>>6��f�"Y+��gY8\�蹗c.a�sǢt�zpBC�NW�'+�爑���AO^{Ў��y9��99�A)v����YM�e�8��q:p�8AK�z���d��B�,h�K�SN��r�4��q/�|��|�ZC������x�ǥ�q�O�̮"����iM��o����6��>,�d��f3Eld��J,��)����S�-��aIR���%����_c���Pİ�%r�pIr����L6cK��Å�xY�26.g	̂RR1�Jk��m
2�IK�J�|ԶId�[�S�L-�So�1-8��
��LS%��uOi�&��-��v���'�M����<W)�̺��ٙ\�l�7CPE�#�Rm,�l����]��=�㵖�}Qh�'H�|����A�R%��Ki|���*Z�Ld�`�jQ�Ḏ!�e�����s�ZgK,�����<<8��p��)�#bu��sN2g3��gFǼpL!
���A��g3��sd��I�6&�؛blM�K�}o�/�o��e�#���c����;gL�1�3=b}���'�M�؝�u��F�9,c�1����xhJ-�0�@�F�DP�&��N ��HI�0���T�Q"�Y"�,�E(ZS+iN�q���my�1�>S��-i4FRͮT��ӇN�C��Îp�h�lqL|jԖ4��*_cki:���8��#�a���q1��)�|�n"T�b�q�1n�HvHL�.�%9�O ��w9�q	�G#��jB��"%�-k[��:f�-�/��vil4�㏣�ʹb�u+�͢�r)��-$��ڜ��q��L�H�dm��岅#%�Z1M|ȗ�m�Zi�i�����|�X}%�J���\K"��TI�h��ЪR��hb7(���g\h�q�>R���C��(Q��R�H�F䠩E4�8[O��%kۊK�L�8�8��ȍI�"9�C��~�����g(��Y"��-��9򒔴Ƌ����t͓����dlO2�#̯b��y�iŜ���I�-N#\1�����J[S��KMS�ijI��d�$��;��*�	K�IKD��S��9)�%N�����0�h&T��>gԎ�cLc��2�e�/gn�y�N�:�T�4p�m�>K�S5(����1��YKki)��c�������6�lm*YT�)��t]8��e6F��M���BV��*�+%�˥Y�2KFp�c�Vq�3���3�JE%QSS��ϝZ�%�4��JL�Өe"�Y�BT��[d�ٷQ��IGҲJ44}-�|���4�F%m���;��{��q�w>>8��>:al��B�(�������MJ>If����%��D�1*�K�*��E��KM%�џ#J�|�H�;1��YQ	Z*\��."T���gާ_%�-�S�u��ckSJc��o���Q�NM8!�p�"�1��m��M��%���ϛi���>S[KS�b��|�ь��gCM0���ɕ����p�Je0g����!Du�>i�R��N4۬|�$�0�M>[M:ƜqM4���%m�a�����!i8D���DzBh�2�e�!�C(�(q�!a��!B<C,���o^�b~<x���C(�Q��D2�e�S�(�Q��!�C(�Q�D3�!�C(�Q���!�C(�Q�D2�e�!�C)�2�B���!�C(�R�(�A�!JQ�D2�e�!�C(�Q�D2�e�!����r��Q�S���u:�N�S���u:�N�S�����u:�N���kZw37RZ�N�S�g����[T���u:�{x��uN�S��L��������oU�qff:�C������uk��:��;��zt�uF��wn�����j�K/�D�}w�:�^wΧT�bN����Sݽ��:��;�S��:�\�ʧ'�N�ծ�T�N�U2:�ݕ^O��S�]ܩԝ�T�d���uc��ھu:���7I��i�_�0����!P�*R�E)DB~�)J"�t��cQ�Ds)�(�p�JiN)�]4���"�!J3YJh�!��(R��N�!��D2��S\u��6����<ӏ1��k�Z[�D&SFQ�!��e�!�F2�2�҈��C(�Q��!�C)���єGE��D2�gSOC(�Qe<2��/�"�)J"~�D2�e�Q�K�<!�C(�e1�i
#�DǙ�
3�!�C(�Q�D2�e�!�C(�Q�D2�e�!�C(�Q�!JQ�!JQ�D2��SHQ�~u2�e�!�C(�Q�Dc)�(�(�Q�D2�e�!���<1�C)�2�"�e���mRM�ݵG6]���w]]T!�!�=�B"�☆SFQ�<�xe�!��MDq!�C(�Q�!
R��1�!N(�ze4e
|�SQ���!�C(�m�vU"N�V;�����{�YO�G�A�1�D2�e�!�C(�Q�D2��8G!�C%4�e�!�C(�Q�D2�e�!�C(�Q�D2�e�!�C(�Q�G�1�C�Q�D2�e�!�C(�Q�D2�e�/̢D2�e�!�C(�Q�HB��!B��!2�e�!�C)4��!��Q�D2�e�!�C(�Q~�4�!3�1�1bD2�e�!�C(�Q�D2�e�!�C(�Q�D2}�B� �A�!JQ�!JQ�D2�e�!�C(�Q�D2��(�Q�D2�u=��L!��)[o�ڜum6i�1-��bT��\ci��Zq���i�!X�xÌ<O��%����9�L���_E2N�������N}vd��wb�����"���w��o,�o�M<W�ޛ�Hp��߱��x��B�cf"�8�(㕷�ۯ7�ov|��r�e�Zd�qHiO�#�-��u�q�:��K�%�M��0�1��r]��U��Jȗb��r���[׷ZÊSF|A����1�m��uM:�Ĩ�Vcƚ|Җ�V��|�lum�,Q�[m�����<�Scڦv�l�|X�Bf�,��8(�Ɣh�2�q�!������/�["G_U���ں�f�4C8���a�0ga�q"`�!�LV�N�.��W�5t=�!c!���F���d�ؙ�`���Dq����fA�M4Gj,AX�`�#Īy�Y:z�^���D�u:�N�6'�>>��~gI�;mĩ��n���bM��g���8�ў<}MLТ�U{�u.�8�����0�Dqǆ F�R�S�:�����)��T:���!<aF�Fi)����4��<q���f0e2�$ĭ�/�n��1��4c � �CL<x���wLZ�l�y���Fq��kuK[�)��ijK��[(���6�t��6��z���9b�1�ַ�%LZ�|���h�!�0F�ǆK\�-��~���ui8�Kq�i��꘦<�cjm�ֵ���q�4�[qN-��[��lm�:���[Z�!���w˯tI��������3�xd�
|q�q��JS��#L0�
"m�_�A��1�[��J�۬i�>uJS1m���M�cJZ�>K�6�0��xb<h�a� �a�߷o+�����/�xB<aL �2���!�C8��)�0GǼ�ǈ`�qD3)HCH#N �A��)�������4��S��ٌuki�{˫��ێ�8��>q��8�8d8�!N��C�SƐ�0���p�SF|hi��0_�zڇ{�%�<�Qg�!��ƔE�!i��h��8��>M),B�4��Z�NfwT�y���S�mjc��R�1��򔡊�$��aGiE�,��4���cjK�Q�%�|���SiY�b.sg�`qCŉu�Z�#�`������ӊq��c��p�>��p�o�g�M4��D��AQ<nM���ӍG�)O�<q���i��q�M��O��e��c�6⏒��0g�|g�C4�� �Q�D2�g��<SM0���F�#4����h���iǈX�3HP�0�B�8�;��a���Ŗh�4�!���Afx�Oid8�!!"�q��4�E8�2�<|q�1~B� if�h3�(�4҆!�3F1���.���(���8���iJ|2�!F3N�3�Vq<uKuJmkZ����S�K��K�qԵ�[cN4�Z�L�u|>mK|���������1�D?�!�ݓ��W������8�M�zc����>4���3����Ŝ#K0��8��"up��JSN4���.w�i
q�q���"���CM8�8�z̾�e[�h�Qq��-1�c�xaF��x��3��3L>���!�
hC�)�p��4��<B�1�4U��@��5YF�fq��AG���_1�[�8Ѵ����4�l����%��:KIjcmN�.����0P�q���؄q�<|N��|P��>�?�i�b����:��Zh�m��n�Hq��k��!iᆞ+�7���Zا��cZ�K��g)��u�G�1�T��1��u�).�g��A��a���4��R�}�%�?�gwaN0��E)�q���ԦR�ckc���q�q���4��6�KO�)KSM(�����YnB����/v:��J��)�ᔤ4Ӎ<1�E<1�B& |"�a��4b�)i���wuVI>Z�h����b�l~s��f���y���/W��!M!�M4�M0fƞǎ=4�C|"���>0�Ba�4d�����gC��y�"�ktѵ�ۊ�]�Q�� �!��(�f�<1�+B!U�.�3�B`�3Ma�>4�DaJ#�q��1}��bu;����w�3�0����cEYc0ԗYFS�8��F�p1��"��B��H�L;�]swۙww"��g�vn�9T �A�bQjS����rc�K��i�c��Yf(�4�:S��v��^��{�iz��V3
iLa�?���G��w^����^SLuKu�6���OC�a��CM(�ح�X�s�Ӑ��۔���G1L��ޔ�R��fe�a��2�3L�x�8�BBBC�!3�0��aHq��
`�h�!���m�'�^���x�Z�=d��mۏ�'�31��u:�On���=�~C��Q��4�M%-4�|�M)n27�i��8���||Q�b1�͙��1��"������'_{�qߢ��
CH#D �"|`�a>�a�M�f�b �x��i��6�i�퓾������wb���~�~�c����*���m����;�����g�cu��|iĴqlc�>Z֠��YB���F�aD!QA�D2�fC �8e��0�Řqa�g��̋^�I,���ݑM�$�Wf��=z���g��{wq����}�㛻������N�S���\���N�W�}����4Êq��(�Q�Ҍb�Q��>4�!#�N8��lu�-�c�����)J����8x�pa�#H"C(�Q�D2�e�!�C(�R�C��t�'���=�����y{$�d�g[��/�xZž{kuϯ��5s�ݹ��{n�']��j󯊭N�$���l�8�X�-JS|�:�Υ���J<"�a���oҊ,���34�a`a=$��x'�ms����%Hwv>��$��T�35+�&홚��Y�RN�]�WUD=��߾iz83O� �8�i�J"�D �x�L<^���K%?/��Q�Ɛ�#8��qDw^nܕ:��K��u�v�U7�N�S����RLK�$�ff6ܽ���!�)S �C!�H`�"xﲓ��m�:3��8c<"��wj�8��$�ٯi���{�S���߷��{���Su$�[�1��Va�!R�D!R�F�p�p�8�)��I�֒n�Rk���4e)�)�}-�3�ͫ2���IN����M���ө������[�PiR�� �q�0��)���eYe~=싗~9C������Fxc�)"��a���2�c8��!�{�}����w�G��8f1ÈB�qJ2�e0��∆��!
Bk�}6߽�{=0��|��Y���,���7��b��)HBA�d!JA�M��x�9xe�����O[��N)�%�����c��Q�"��3�(��<"��<2��!��l�R���C�|��r4ԧ쿴p��Kn���9�4c8�2�ٝ͏��c�aAF�pB�Q�4���ܞS;��η�-8c4�� �8C,e�YC8��`�[m.�*'���xӉ|�m��IijSLi$�c�R��Di�!~���3/d�r9s}Sם}��/]J���2ezIs�}{��QC �(,�K�D6��V���aiK�m�:��7��b]�>��gN��y�Mn���1���m�0�i@�!"�i��@e�b��p� q��!FiFf,c!-�y�W{�ʵ�=uT����yTj(��K0��Q�q�8��DS�Q�G��֛u�)Jq�>iImJm��۬<1c0ў8�8�4�)D2�g�꘼��N�S��~�w2H�R/>���[�7�<)1Q���D2�e�#�8�(�<#O�]]U[y�*�%����.��%������8��QC!�c4�M4�>q��K�6��M����]J�ih�`��ۖ�J�I�snfe8��2��!�C��CN�Jp�2��_�y{������.���!�#ǈi�)<B�qJ<`�qM�͑$ݒ]��M�fH����i��!�C)�d>0���4ӎ
S^{x�nW&#Fq�PQ���!c<!�aN(�X�n��n'HBZ[�)�����:ө|�V�ZQ���Gƌ��SHQ��o��#� �!��4f�q�r��x���q�%�V��w>���w�R�Oc<Q8�{ٔ��D`�3(�X�p�(��8d)>��Rv�jK[Nfek��[Ku�|ť�'��v��B��"�Xi]��U�!11����D �Q2�)Qz�c*:S��lR�ƛm.���m%���`B����2BBh�4������/H�N�S���u:���q��B��0�8�0�p�!Ja�q� �)�(�1�0�8��4��4�e!Ed4e�0�8�<xd�!���i����G3�1�C �A� �BF�i3�#J"C(�Bq�)1��)`τ3M��2�D2�eǾ_x���<a�8b8�2��)DB�)DBg8h�g#�2�2�B��BA��<qiBe!
R��!C<1���Ϗ�!�a�a�B��FC�C��!��<Un��1�3M�������]im���|�]mIm��|��-��y�~�-��S�|��)O�ی|�1�����)��ь�N4��N)�RS�i�'����qo��̞����FoV�u�1�b�2�fC � �B!��/vΊD�ߩ/�i�X�Ĵ┧q�8�V�e�;���x�ɘh�R�^<R������T�uJ�N��lS;�ݼ�'���u:�N���T������uff:�N�Vfc���bo����D�u:�N�S�[T�{������O�=}���UJ����I
�k��*��'R>�ϵ���E��{�iI�T^�=Qo"W�J�I����:�M����8�'�Q}Q��|R����CQz{�� ��e��ѵ[V5ja�3ʬ�=��{D쏨p9)�Ou#�8G�+����_h_b]+�䗕��	_B���=�HrW���O�N���aL�|P\����ӆffq&X��S����߮���c���$>�-��a��L��Ҵhi�a���bb�Nz�&Z�S�({�4L!�ܻ�B�W�)�h�3*��L5=�|�EԎT��ʞ���/uQ�{G�"��^��K�H/P��_5TuGЩ�_iK�U�<ʎI�Hw��@?���+����O~?ӕ�Ts*+%DUU& ���v�K%6�e�I6��9q�������G3���r���Y���[�U333����:8���3z��ʭ{v�%s7feӭ�ʞ���r�nr���fG2��=ėX�G9[���9y�]��ꈍ���*�}Jȇ#����9���ͻ����+���L���W"yx����"++�͚��DY�#7�#��(�"BU�B
"j�*��+.fTiݪ�����r�\��誚�$��Λ]u���1�vD��)L%����LL��7�R9l��\����"=�TA`��
��$�1�D��o)�R,DHg29ʈ�G*3��r�y��GÌC�6�����x�.�"���E�W��Uw"H
D}�>i7��S�-2��YQ����9\�ns$ ��y
��#�qQD�S{�4�ƪ�F��V-F�.�"2!�#Jƕ	A�����d=���>�\F���r�����*X���(�٤��Qƺ��nK����U3Ke����%ԟ6���Ԏ��5���L��6�-�o����q��q1��ƻ�)�^[Lf%���I�����>��׉І�v�,q2J�ib)��:�{T|������~���U�$dX�ʼ��z�1�1��&elZη՚k��k���R���R��1��ju��Ls��A�,�_,�Z�q����|Ī��e�2Ru�-Kru�Yƺ�i����[kUF�KH�]I��Y����8�ͺ����*��1j�qά�����I��f4�Ѽ�h����o"��+2��M��q���5�A�â��2�I�޼���'�f.Vg�uq�ţR�N:�̄��bm)���KR5�V|�rq���*:�8�ƔĲ�)��v��ilDAq����㫆����J�+��/�L!	u��~⑝yg��j;u�Z�Z�nZi�|Tu(�*;��_eF��V�#��r�s,������F��u�\1.;"_}��!�A	`�z�-���l���ѹi'}g���C��1av#0��@Cta�Tu']}f:��4���&��2qo�>kk�����F�䭉h�Ɠ�R��^�'�R>k�n��{ߦ/�9_��>fT�W�˙\�ʬ�U��ٙ��U<ʦv	 �؉��"@�S��ٝ�tEr�j�2��,\�'y=�ˢ�Yʥ��1v!.�n�������A%��JB	f���Rm:�����,İ�'+3-�|���JX�M�2&�"���v��2ؤ�\WW9�ל�Y��re&14�/N;H���gT�co�i$��>��&}��{�z�Y��bqM#��M�ݜN��q���R�E|���Ҷ)}՟|��N�����_%-7ڪ�f����K�N�s�}R8�vi.��*|�I,M�Y�8�Vm�k�2xꍶ��i+i���V/H�]��Y��TX�TLhB�Sc4��B��تS�u��g�|�q��Ӵڟ��2z*=]��d�Fm�Q����W��r6���8�*�*�b�9ީו�7���e����]�{s)5!ۋ�B�F.%����7%Zh���J��K1�-u��K1St�u�,�c(�^Y���}|�Z���5����7<uO�8��G��g�j=���Zض-)�rѭ�u�8��T�[w�Z�Ym1����r��|��WR����k}���ؘ�R�k�����c�1q��Y)b�RR��!y�8qJbz�{>�v��E��u*|�
��)�6D��Jct�ga<��>�=��g[�Г]yp�ɗ�[�.�HKv��~>���W��N���d��p1j�̸s���.�t���s}}tgT�cn%��;Җ�F4^�Ωg�8��Tq���M���f)+[��՛n��u�-KrӚm=]+-�kM1M7�W�3)XZX�!���2��ޫ���-�T|�#%��gVd'N;iL\˙��U'��1��Z����}՟7C8�ε]I��:�q�1��\N����7��g\GrὨ���J�w�Ŝo�>Lo�&"B"�WVu�FGcN��R�I�)Y-4u�u(�O�Kr_\1.���)�%�K"8�S�8�$��k�D0��%�;Ll|�Ň#�H0�}<Q��z���ǝI��dLlR8���"��b�:��|��WR�Dy�l��-SK�ؕ*��2pמY�|��:�r�XĴu�I�Z�Z��Gꏛ�g[��uf���JX�R��Ț���K�=h�.I~yc�gy�C��tt����(�������fh�Eg2��Y�Q��Q%V���Ȏr9=ٙ�r�3l�FU��L���/@FXb��ĔxgWE6Ԃmq��y ��0��j0�J%Q����N7����v�o��>��<�8��8��٦��'JV��u'��Y�3*{[Jr9I�=ʵ�sWuJclR���щ�mG����)�W̌M$�U1K��qL���1�S�:���J:�v��E�R�}���i6�)��N�|�r�N3�4�{+�V�RR��ًGufۡ�[��WRcm��u���KU��h��y�F�mfuO&8�%ם�oS�8c,b�S�k:ߖr.��KLZe�ė�wi����$7b������#�g[�wm��T�fi��!�%/XxVN�)�)�TB��*���ȫ}Q�Dn��ʞ�J�V{R�9��5�QS#9b�'���s5��Ȍ�T�׽�vfk�R�FgFN)Rb���Ty'ϛ�y�E�՚�G_2�Wk[ť0������3�,�|�����qx�[Lf%���_P���:�GRu����[�U���ԩk�=%�<����ï9hԼ��.�uO�k1mN�Z8��H��ڕ+c#U�2֥'D�H=�JI
aO������u��]'kS�Wq&dZ�J�N�0�NKn�C���N��H����S���7_Gb���Ʈ4�#�u�.2�,�z�#���m��LR�1���lZ8�m��Qֺg��a<:*�xf��``q�u0��-�|ufBt�6�**)kJN9՜u�����W2�Q�IC�Bt��(h��1��O~Ɵ7g��ѣ��Ɣ���t0�Ѥ0Wț����D���k8�:�q�.ڎ�1+U�/�F����}'ugZ�Ј%����˫^iKZ�-/P�Z>kk�8��v��pa��p��$��!E�KJ8�҉te�����.�2Ι��c��7�/�#� �((3�Za�-�Bw�^��A)	E\�s���t�5�T�]:�WR��)����B�6�.�f`r��0N�3{���Kǃ'8�3Y�Z'���7�S\��Srmj��n[�˅�+.���Ǐ:v��=+8�3�ӧJ�<zt�tgҽEåNՕ���>B�`JB�%��\!��+2�8��cY�u�v�E��H�DĢƩ,R��${�>Ws�9�W���3��Ln��;2̙�+�&c�Yf\gcdՑ�8Y���g3<6��Jec)"i*XT��4~uե�q�f�efG*##�����������!&�i�S:I2���i��$�$���M��M7*9�{"�WG"�####:2�'�27���#""1YQ��u����Έ�F�kUU������������3�U����ޯUC�]gh�4�kI������%0�k�'Qb�Jb�H�Ф�ے�ɡ��W�����sg3����r����G+y����s*�\��QY���9=��G2�9L���;����2;9ʮ1���dr.2�Jmإ�DA�
�R/c��˙�����r=�\����]r��_7*�fb7�QTEC�Lbc2Klh�y
B��aL"���:&fdD��Ufk۷o]Y���Y��TN�w���+�x���$�řrL���!JR���nV��(��0V�r����	B:^����4,�R˲���U�VSpLݓ\$��9P˧Fe��eU�Es��1��!L���Dz-�q�gJ�V��:vEr���smk��Fs��^�S�ψ��<<)H�( �Y�"iw����ٙ}]�"'�:�K���+9ɼ�neR���ʊ�e�fT9YLdT����̤r�����UqKΞ��c+:�ͮ�;e�u�7?NJyR}�RO�.���z���==�"�Q���G���&Tj>p��g�q�QƓ2y���;i3-�>=2��%:��2ֵ��T�AI�%4�����L�g�n:�4����~b��&����'��9Į���h�b[W����I������ԙ�f}���ӎ��E�drz܋��Rs��3H�ʏH���Bt�b��fO�\?2v�f^ߟ;��_{�ϕ�>Z�fDd��$Fuu�;u۞T�Q�=�q������O]:o�QƩ�>����Rg�&i3��NQ������h�Pժ'k��W�hm0����㎟�i3S���T��'箝3Q�L������������3�3ʷN����8�L�fO�|~b��'�g�Iƣ2y���ڦj>�u~w'<��iLL[Q�ҬL!�L���NQ�L�߷/l���ߟ�|����OO�Q�Y�n���sUDUs3�W\���frJ�L�]�r��ݱ*/��d��6�N��K�ik\kη9[;5V��r0��C����x�JS=�r��'*��lr�seeFZ ���q
&���~��Q�?�e�11��ܭ��\\j"4�[��tf��~����5Z����U���ŕQU�wF�K�])+dbqj^���Y�tq(#�nH3����UE3H����RB��n'����eHȧ����'��:��Q�L�����'mFi=q�Ԝi3'_�S��%(ڞ�s"��DD�Zii�5���L�����;jf����S53O��=c��jo�\u���>|�W1�L)�JV�{�Ra��)O�>�N1f>{q�ڙ���~g53/�����L׷��|1�Zi��k)�1(Ja��Ɇ$�ɽ����N1f�_�z]�3S�ե	L���)��6�m�6��=;�zd�M��2q���R��"���Oً�Jc1&Qp�[R��dA`��b���}����L���2q��y�8���7��j�Uz�"J֥�j�UyU=�2�����or)�f{���2��.{{+&�cu,+�ڡH�Э�u7`� �t��D���0CM��㱎F��G)nv,+6�*����3S2��Ϝ;jf�z�{jq�4�럚vř7��;�>�����m0�m�j[i1	jg�κj��S4���ܻd�B|���E%	L<�?&�%/�[�b���J��1jN!I"R}�?4���׶q3S2��ϼ;jf�z�~d�Go��돏�z����z�<^�����8��N53/���.ڙ����ꙩ�u�na��Jb|�?-Nl�Ҟw�}��d�?=���lY��)����~����ԎFvUDoevTYKUҥ8�bո�!I"Rk�m&&!)�y���R�:�__�Ȕ�=	�i�z/�'A4$�,-0�LK؞�N��~(t�;��Ɲ�fO��u�8��&yۈġ)��>�KUy��j�lv���fL���휅�����{d�c��?2�����H~� �A���U;���Ji�6jJ������)(JQ�.ڙ�����N2gן���䝺�M�kLb���d��"""���)�_R�2���be3���������
�0B��B��y	�'�S�̍Y�9س�et�B���?>�����>^�h(��o1��Y.1-b�/4�b�ľޕ
��DZ�3��_������S)��^&S/7K��m���;�ň��$%��?��x�q����QO?��O����|�-Ji�ST�O^z�2�}?.�-�4�q3��p�F�-���08����W��ﾒ�.��~�K񦾡�D�eKkl֧���~v�fz㹓3>n�2��"���S��n*�ֱI��zT�����4\a�?����A `�!aa5+�W�J\N7�����Zx�i$E�t����J2A��U�a/%�"b	LR�e���/��ZIC���H�Ji/��n҇���YH��Y�+>�cKƳ�t��ri,��ʙ��^g�B������mF���zU>�ŋ���4_��~9W��~4G�9����X�a�/���i%�8����o2����(ژ�Vc��c{�U�����Z�)�3&�A��97T؝����^��CNr�����}y��X�EW'���fՑ&�mɜC-���+�Nra�gb�E�,�	h��Ȍ��g**b*u�Ͽ9���)|��U�ͷM-�Z��9_����Q��!0��uA�	qb�)M|�~?_J���fg�_�S���E)�����%i����jB��ŦQ�E~�?�H�I~?n�^7��,!�?|���r�2]�:%%����.�K���+�t��~+�K�£J8,�
�.��/~eL��neUO�����n.������37m7����7��󿗓3���R�'{�|�~6_]����R_.,���1"�������q߉�E���&�iLb��C_G�����|]%��3����#�+�Hg����~��j����r�9���ӗ��J��2�z��3"1���y-%��F,�
8��]YYX�d�s��gW�1�PЈ�5M.*�MYM,X�b*Ш�E��I#W��ZV�3=}�������S���-x�kM� �����8_����_�⻕3/>������W��v����$K��g��Zo���1~%���\��<q�SWl�j����Ȉ���*g�G�S:��əB	�u�T�Ýw��XɔYX`�đ��4�,?I܇W"�z�W�ڪ���1j�DGWZ��8�2�g�����g��Hi�����%����(K��K�C���'�ƪ�9\eL�����d��Q���M�t�r3z�XŴos3=s���&�$�����EO���<�6N>��ϳ���<�/��xa_"�����Sτ�w�g�=���������}=B��7�X}+G�L~\v�g�/������0�""*�?+�S�+�Iuikʬ��Z������c�<O�)
&�R���rFNm}ɞڢ���?u�T����ʙ��*�u~���V�ݷ%o}��D)s����������xX{�_��?�_���r���W���__��h��?��47x�dO�*����B�ȅ̸�\��}�̙����}K�4޺(���Q%H� f$��SJx�q��"#�D\C&|�5�3���ɟ�}q\�SXի����~��ʙ�7���ϞWr�Q	y�\�4y�q�k�������^w3?�~k[[�ȋ���I����OečɌ&�57����~=EO��U�+�s��<��NKi����L�	��y��t��~�/���'��Y��.�^'��_���*�rY
�3�!SG���>Zd.�^?e�����TD'۪K��qq�T�Zi-\ϕߋi(-:�>>^5���D���D{�5�ͷM-�Z���+̩��_w{l��ζį�̚Z��FG�"Yq\K2ef-�`�&Vɳ.&��g��*�2�DU�%�������eDo\�����2�:b ����LC	G��J�vC'�gr{�\̑{#$R�eT�b�z��5 �ѷPI4�Z���b¹*5j����EDu��Ti#�������+;K���{��~.�����E��-�X0Ē����~����!����Jc=�j��s��ppz??���Ix_������C�a��ۣ���;3UwǞG���R_J�!���_f��=O����O���/�D3��e�XU<���o�� ����w3?���ʙ�������\�ێ~%����֙M�fg�گ���9_����K�����z�qg�<1�y����8�~?���W]���5��3$C��~~sL��'��F/vޛ�Җ٭L�������ҹ�E���޹i�r9YUk��#HA��R�G�q��w��y$������m%҇�Gp�e��i�M�'��(J)D��].R%IR�R����J�4R"I}��Y��i_�����Uܛ�4�`Huz�ch�@O^{�켨�/��Ec����Ll@�����ۖnGޡ8.�l;�����<�bZ���O�/��s�t=Nև4$��H�$�L[m��	%*i�J�$K|��m�Onױ�c���p��ǵ8z]�2e2�q�v���
%(�%�����
	%����d�|Q�K"�%bq2��ܔ.�4��E�Y3�w�o}�^�,�阮œ)ǧ�L��ffq<=>(I
a>>|J�$���S���1L]��,�-��1�c�1�m�Y�I)�f�ku��VZ��r*fFf1q�'B��Ǽ<0��[{ܬ��ffs#�U�3���Zյ�gLW;2��G39����WM�2%X�t�G%v�$�w���ȅa�^LTJS�����	�UV���r�!��er�+�=��fU㚯�2�UsHA)K ��b��%d�	�b)��Pv�(�5hbv��7cj�L%�!D�D��T���)aH��B�G<��qu�ih��k}9��s��F�UgW���v㙝$�Wο4����ޓW#{#%�٣�Q��fr$ON�H،�Mk�̅g*�8����f�Ff8����LN��K�v^����G��Q��TuHq>~%}����U� �K���{�ߤ�1�&Ԇ1��&�C��H�+���9Ȋ�U�}/%/%ҕ�nJP�)v�� ����n�Nrr�*�-s�}��x��3/�9حHJ\���w��wK��+��+��=�/���$!�3/'�ƒ�W��v�7W�eȗ���, IiQqt�1~%������q�Q��b1�ݕ�%��t��D�>�x����_�����|��X��,��JQ$}��ɤ��]�=y�2g�b^W'�*x��]�Rj�X��HxSe�>+?��=���*���u�쎋b���dfG�p��y��fgn�S?������~h$���0��	u,JC����F-l3s3�-�T�έܩ�)�Uߋ���ϣ���y
m�q�RO��g�,���eE!á&:�u�o頻�u��jk���ބ��ip^�����1��<8;f:��s�h�/�1Y��xX��0�@�ٙq�_��v{ߗS?+~e��^r��L��_����j��,EF��s���M.�	x��]L�廕;�Q��%�bo�+S("w���3���ə��d�␉J"!M����6�q�uk��v��k��3�_��wuRL��X�g1:"�lB����v�Z���W�Iq���^fL�1צ\��F��4�Zj3JCsH���(���A�p� ���)�ޗ��S�E�C�U���?Ӏ����`YX�[o��}����罔�5jn[���3S3/����DD�$�$%s=Wz˙����L���~eO�\/��k�-������2gy���{c�G)�T�э��D�e�US[#bl���3�F�����|���鹟4����7�o5+cx�����L�U�}��M����w������:��%$�����p�ŉ�'�	�xB�����}ǂ'�2ZB	C������\0���p��@��b�g�|̙�y��?6���f������E6���$�h��Ņ1��?�x_S:���Ƒ�����d���S���.5j�4�U�����gjs�����/&gϮ-L�Җ�z���Ʊ�mlkS?u~NL�\[�_�!U�Q۩�~~fL�/����k4���-I��Q	A�^�̩�w������8���%|�UT���K#�ʪ̮�OffH̨�ET�{z{���"��Z"���ٜ�Oh���9U�މ��E�MỶ���/�&�i	��p��:�v���0�݃0��U���.�9��ت�ecZ�u��#��!�_�.x�򝊗[�2R��7i^�g�3?�G���_G镜��"9�ш�&�qK���)���>�����{1�|��2�ϒ�6�m[�U']�%0�C���XSc;o2��~6R���_�?��-$��SK0��౎2!�!(�/{�}��%��v���z�������}�~5D����7x���O�/�w�}?+����yǺ�c-��6�-�ҽ�fK�U�����^(��m|�x�ô�B�gv/���b���>~6W��~'�a$�옄/)i^z�DŰ�֐��8���幕3/'�S�%�)���B%M-Sv��Tb�9͔�窯HottZDU�]��\�Ob�9rh�3�e�츪����bW,rZr���"9\ީo�l��,(^�1��������_��5_��칙wʴD3�y��u�~qL)�)����<��=�.x�}��U~���I~?i~0ݶ_��#(�e���~�/�׳g�����?�U�)�̹����-4��2t�4�d�C��6W�e��<���;����Y��CE;#0ȈYfb_��K����ޮR�.JoF�䵓�}z��1�_����ҩ�~X��/�G�~'�����Hn�|(��5).i����/�!<)⿈~>�s���^o�������y��U�U�q�D�~<�����kM2�f|��3=y�g�B��+�*�a<��/�*�/��=����q
���2�e�����=?.�y�R�-����Ŋ�<�����^ミ��������"m�c�xy��?1��?=��D_dF�"�W:5��b�N��6)�o8 �G��b�����4�ݺ(��DD0,��~����U^J�����ws����o2fz���AS3̩֫ۯYSNd��b��j53=y}��B�EO]Z�g�ϱ�3/��u>i��q<J2^!؉d�x�1������|��*�.e���gO7�3��<ť�'�	�y��r�'��>^�>~_�S?����6�����k��R��J�������Ŧ!d�I�	��/f�nd��șQ~��Fܮ����������g����k�TjӼ�|��7�2���o�<�S	��?6W�=�U�y?/����ע[}ꪊ^���z��<�� w�����ҫ�y�������=	����7��1(�W���锑�GI~+?��^+�Xa~��(��'���TOYN����W���e�^o��k2ڙa�3���JC�
z!km�\�B2*�fT�"��US���d9R���ܾ��c;��e���8�L�\��O�9��.��#+9.dIs���1��Lf��;	;2���gN�;D5G2g*+3ds�9{{+2�Վd{9&Oi�Ȉ�98@o���d��K��c,��]�IO��t���R����|��sfE[�E7����cG��$�㝤���t�h��,��)���Z��LA1hi	:���Oa=x�I�j�����~��S�W��������$�C�(�/�s�@���]���~_�Tϕ�7� H�T����c-���SM�zܪ~�|/�E�OᪿOs��=��|�^��N����!=y�əڜ]L���3%��q���8ޭ��xz|���~���~�Q��!���L�oV���Ws�������^v�32�v��ί̩y��q,[Ξ;�_j�|�m�c�����C�C)W&���ӊ��%͙}�2���]�es����79=�U�1��L�K����l�؉�>��u:�DF��ef"�V��F��W9�2�<��M���W��~4_G��_�����'᫆���1J���m�[��y>��<pU���l��U�.C�|����0��oC+��/��J�x�ô������!������HB�/�/pq������?���9�DEo��2g���)�&׬^��SJ����������	/a(��PLcXY�!&M�JA�}�O���Ix�1� #���Fa��YcH��JE!�&�Î��D<���_V�{W��z���_z/�?����eOv��1-[&ex�ERuS?y�g���Vq�\�[��ja�ˎp�2�q�ΔgC���3���'H�J��#�����m��~o��}m�>��I�(B�Q���˫^nm�f崷��?���G�����O��/U����{��eȬ�իL[Kf�a��"E9o��}��ؾ��������>�������A�)�/�*~�%V��8�	H�2�dfG�33����]�t�^*6"�%��>���Z�f?������Tә-^�ҍM�)lU%��aS�Jn�<W���4_d�M�Ϛ���#&gʏ]O[m�+���%�y�^��O�C��|��U>�%W}/�G����C�R��,�̯מ���qqsz��R�)L��T��]uӥ�,e�e��Zp�&������0���[��Sk�$�]��9��v�̲ə1�\Na�8�cY���x�S1�3�e\2�N:x�;v�1l�j��e���N2��3f3-t���Ⱥ�]<:t��(i��&4҂T�#g����#�eTs#3����gfeFFFFFCD�12M4�u�K�\�m���f�M5��-f�t'nB�ٜ���YUё�Ј����������]���FFFDDoE�H��FFFFFtr####""2�Q�=�b��"b��f�ј��'ozk�3#�YJ�T�f���D#��L�q�hXN�Y�b2�b���QÙ�S�ٜ�o[s���d���3*-r����Dd[�U��*3��c9۽ݐ��E�U^V���3{���EeTUʎTq�c�ȨG��;,q�l碣��XMɭ��v-D��"���T_V�5�+�UN^��rzd�۪��F��̎ub��vFr9;�����!iD�1���D!ԍ����\�m^�y�ܷk�mʨ�dr���N����UFTU�κٮڐ�y-)����L&1�D�y�TDwTkwX�6e;,����*��S�!
���V'%�&)La):��B�NFEX����K��UG"%�fD9�w3*��er�z�U5��{+##:��s�����s�䞬��5D�G'#�}�ۼ��ܨ�U+*u�9���Ҳ�Q���s*�+����FFs�����Ez"��doi�C3e�m�ښ�c��y��u;�RN�^��A��Q}�v��T��E�J�����%�,!�O�dEJ���a)�x�	���b��}6W��R�wp/��>j��:�|��R4O
xC̾��������">�B��BI�am��1���|?���W*��g=��UTR�m7��L�m�.YiJ��^1mB�i{�ϔ��g毉ə�ߐC""3���ʝ����t!��%2���?j���X�י�3ז�D&q���K�ov�]���$đ��M%f���Q�t���d�[|�K�5l�Z��S5R�������=���G��W��e��p���t]1r���d���"@��<$��.�fnEV�W"�EnUVr9�C�&�4����ȍ)hn����\Ԝ�O{����v��2�"����+Hѫs;А�H"6��\�"����\X#8�a/Z���=�Y��r�b�/^ߏx|Q���5å�u�Ō�L�H���J��߈ZxS1�!�-�XMŘa,[�^i�z����SIx�9t�����hE<��1����ʬ䙊���{2�5����V���Ig��.���cK��?qev[�
�0�$�#���
J���%��ƒ^?�/#h�>�ǖVS�xR����~h��|,N�_Õ�O�:XA��G+>fU�"^?iL��>˙�g˩��y�2����X3�S˿�$�~?;Ix��B�1
���H,l4`��cET7��>�K��K����%Vܵ½31QP&	6������uݪ2�+$eʈ��>���{�rUG�r�i"9�c �KH���V�IJa�Pn [�'cB�r�b�2��k��ȎW:�fy�Ӹ���~��C�U�������eLϟ����_=o�[3X��T�M����w����|)U�ە��ʴAԅOߢ\s�)W��M)��z���~]L�վK�?[^W���x��մ�iM+DD:����gU������5Ke�3�^�{�y���!�!z��c	�"��ec-�Z��DBqˏ�qo5O'����R["���QS�ұ�r�^ERt���[o��^r����v<��ה�/R�鎼���WA1[��I�bW̓1����D�|uϩi��ן\""Ƀo����I��R�����r��ӎ_���_�y��>n�g�5����SE��
B��5�u/?>����'u��4�KX�1�E����~�B���ִ�1+��p�Fn2WdY�VY�h����ߖ��|��߭��y+��)�*�|�8��V�Ls*��6i�<��|\i�,�]W�����R��)��\���5ź�}��'o���yx�SSX�-���~���ֈ���y[�{��\��Z�M-�5�y�ۮ�o�ˌ~�������.Xձ�i�y�-箊Ƣ��L+*�8���ŷ+�{*VS���G���u.����li��̊S5�s&D�K���z�*�r��-G�W��8�u^~Q���m�g�_��YlS2�ڶF߿-���u��Ω��*bf"���6������j�YLӿ��7����-;巧i^>;t������"�[E�������?~Z�����IS�E[��_eEZ�WVgr�#u�1�cA)<��DD���4�Ѫ{�s�U���Y�eVVM��5Ȫɗ���J�^�mȽS�qͬ�^ʑ9�39��ќ�%$�[�at�����!V�+�2-�y4H9_��7��]%W�dJ�c�)�/-���)$v��Jj%/B���x��%�O��̢��ݸ���������կ��|�>|��Bf��/Z��G��fqM���Z���t���1X��4�4y.�F�qg[��N����iv��I��dVcH�\8�I�|�:���^|�q,cM1��z�i�^Z1���_yG_yf�K뿞ĭr�.��RQ����yR�IVf����.l�gY���܌��[�"9�:������n��l�1�~ߤs�$�~��esj��Ei��ܑ8�y���VWI/9=�̓�j��u��"���5�X���tdg5s[4��=��RW#.C)+cg�yh�\7�<�c�Y��m��ʼ[M4�l:�k��Q�޳}Sɍ��ϒ�Milұji�y�=&�qfy��9g���J�5�����5��K(��,�!��i�������^�U��G�㟅L��qz�{9��H�M�H�K�'\s���S�i�,���+�k�Ro�e.��.�U	c�)L�b�<��4��1�.K�)��q*�̍-Zb�[���?3ļ[X�`�Oh[��:��|ߖy�w�<Ʋ�֖��[���f|����O���>����߭sNd��[ZJ����F���u^H�oY�ͼ��x�iy,ĵ�s�)I�%N��8�Ur�o+t���J��3&�8�d�>Y�yf�w��Y�����BxB�\"h98�<��juz�:��c\Y��Z:��6ӿ<]f-tҪu�-���=p��N��y\�o{�ŭS��-ZRT��壍9l�"">�OT�M=���%���1x��le������m�7�<�4�{�Jf�S�i�h����ݺy1�)���ZT�.q[3s����ڷ�)������6��眳M�ꗒ�Yjj.���Q)�	ʣ�#睩�0z{�6��G_yq��u���^1���Wz�f�uO$���y�rQ���oNҼqLUZ�Kza瞸s�m&;�}�m��IU�L�S? �����f��䶈>|��'�U$���̨�UVb��=s�����E_H�u�^9^ދ�5b9=�ܪ�w�����9ʎ�"�4N����"�O"�U�q��J]]q<�n1[�8����B�q�ݽj��ؐ�1�bT���^g�� ��,�8��ĲՔ�%LkR��z��7�>��|���Ӝ�λz!;�eM�*a)S+h�>��ѷY�����m/�|�ilĵM.*�M�Q8���ZYX�1���h��jz��u���iv��M+"��VcG\��"�.���m������~~q\K�Li���1��ה�kk�~�����~Y��]/��%k�ZV̖���?Y��-o˄y�91��w֜�34��I�~S�?�1��ăD�ފB&�%1�kioX�d)lb���n~qH�~Y�co���e��#\�Q�E	w7G4��;��L��2��Y�]3��u)�E�6C�%:3�6K:�����1��gUvdffg28�]���s���i&�La�r'��Y�������fg9UM�ٙ29�}T���s33���fg9�U\�)���)]���D�m��a$��=���9��dYH˧*#Dsg"�R�T�V-G:OT�;��1��R��Y�*�25r���W.s�rUXF�#-s���3W�ʎDUv&N��Y��+3�l�����:#��ʧ��buvD�%kff�Ґ�J��Q�elr$
GzXV[;q��
`��-Jb�dT����KfuVOtב�R��Ha�J% T�*29{�����2Fr#\�{+7�zʍ�]s#�Q�*�)�̪���n1JCM���ӎ�w~8�|����U��p��ww|��Ꮵ>�%4�!H����R�d̩��e��B��a���Q�u1�4����s�Y��^�TuzTT_k�y�۽5"���r/�t�������>}嚞%Ğ��7זj5x��4�iX�4����|r��I眷�DK�ߥ�,���f-u�i{��%��y�嚞���Ym*�%�z����ߘ��ş���a���dmוȵ�it�KKƏ��򜊉���Ds{*7l�D�OFnmȬ���Fe�����F���K�SM��%U9�����mLa��&#�c$)�S���%�}�:��GZ��5��<Ʃ�b�i��y9�Yh�%�"b4�Y�i9���՜s���kF��-j��&VgqWY�C2���2�2ɖ�V�%�=������S�cͽk�s%�e����Լ�s�2z��u�ǟ<��q,���j�#}yf�S釟zε�m�1f��^/U����GU����'Y��u:���F�����X�R���6�ܣ���m��ś*�P�����GfWr�������8��Fu�yO�4��ũWY�L�[I�ϼ��DD�|���}�F{��z%���L^4�1�)�:�d�������0��-Jq���\W0���cڳmyf�z9̥3I��LZ�Ə�~~[�������~o�Ͷ�b����u��ֱ���gT�~|��#��2B��!�1��C��c
�)�|��k�d��G�|��RX����--�״�Jg3�GU��Ֆݧ��~��������a�޳��^*�K��4������w�:��S!��Wze%ja��)}�:��Fy���_�ڲ��Զ��<��\Z:ߖ`���R�Z�R��.�����fd���Vr��Q6^l�9�3{l��%5c9QZ�E3���c�s:)���rDD�&G9��'��Y������*��u�gk&��%_Ef\�����erd��=��OEVs�vFDڲWqߒ��r���q�m/18�4�Լ�Zɘ�y%�/�I,RXM�2�d��b��s�8jvڑ׹f�K��8�M����kzшe����IJct�m��}��g>|��ϿY��Y���b�i�*5��SP�\�o�y��}yf7T�{�)l�%�d�Ja׽f�|�g�Y�<�i���kfimJZi8y�y&���Է��i�c��Syjc�/H�^Yח�Ҙ����E�34����[��+gR�{�^I������q����TҙO�?;�����R�=�KL8��%��r��W^"ڨ^s9������g9�V�{Vn�Mж�:^�LRs��/N��j�}���6�y�<��̌�uYq7�%�]�W�S�<�����>�����h��[�ZT�b�S��m��G_yfOR�X�Ϗ,����e�::���D��Dy�Y��Ϣ�I^2�K:��ߔg|�� y��6���T�����b�[F��~IN�+%eŮ�,J��4����/�����9'���kk�y�SU�ZL�MFv*&6�pLb�����g)��y���o�i���M9��2���h���4�Af��̞��s�1��-q\J�iX�V�G�yfm��y�Y���X�n��Y����E�s�Fo�:��Q��Y�v���bW�Jqjj0�ݳ�b�KKIw�2�#�3=)j��K�9�j�),��q��3�.���V��a�Ὸ���+E)Rw�zk�ŧg��'r���-�,�e/>�ʌcJim4��|��!��.$��,��i���2��-I[J�ѿ<��q��`�L�M���.qbˊ�e�e�fc1��=IWo�q�'^zͶ�*�q�b�#"��4~DK�ߖo�q'�~Y�����{�]J��צ�w��~v��Ny+�iL�\��U�W=[�3.�����e���mˈ�^�|�c*٦�;��Y�f���d�����:���rѝ���K!��UqzK1*a���N9�:��G���m;y.Z�1��cL��s�i�q'^}p�Ϭ��M�8ɶ���Z�h�T�O�qp��y-%��H�9Y%Mwm��s+2�)Ⱥ+FFr���9ݽ��t�����I�		��CLa-H&5
�X��0��0�K�נ��٫��.K�ki��4�1H���9!����E[Y��LA1p"$ �q���{?�8�+�K���T̊�#ϼ�V�J��L���ƎE�we_*�&�lJY]}�u'�rη���8ʯ�>w/�_"���>f�neD�/2�S�u/;Fo��<�B(�y�.���i�jի��M#�ݳm���k�<�G��m������I��yhӎ\:��Q���m��~\�K1�4�î�p�Z:��u�>��mǊ�KJf������Iךjn�J��FaJJYt�ܱ�^�U%�[�;�Nqh�Ϭ�ˍZV�b��o'"��̬��*#�ܝW�{۔��d�r�r9�]̮nZ��К�j$�JI �i�*a"%-/bN� �N�&)�F=��Wח+����1;1���)��߼�>S�oˇ�r�{�ǖ[K\��ɝyNI�[Y֪<��}f�n��E��˖\U����Éq�זgT�[o�K����)ZJX����zэ�μ���^Y֛���5MV4�1�5�<�l�.��U�rs"DFG5WTU1S���L�1,��qm��R��cOS�*s%��Ԥ�V�I�Z�d�*m6�E�h�T�M9���9h��Y��yk��T�J�b�z<��}���" �\J<�,��y-4۶�i-E�YQz:���}�,μ�u�,��<r5l�ijf?%��Y�T쟚���_�{�q+U�&�i�[I�>�I���ծ��TMQ��S�%N�^U�޴��:�&6����3��r&��Nb�_gy���Ffh��4���O�R:��u�7-4�=̥3KRV�[M}��q��k�y'^n�6�*�qME��yյ��yf|�g���ġ�B�S�zs������E8�+чe�7\G16}�g9���u���8���uNVb�[�#���O�}�Li��;SK��Ѝ�kI���6��q��gNpvx�xFQ���L�pYc�g�����K�x��d��e2�&���x����s�=���s�bc��fbt�ヴ�)�	��YBIL�b�c�0ȓ9�fVTC����,�U���M4ӛ�6�[u�[$�t�i�M�mt�UUG2UEG-r���22222.UDU��3222"#/9�=4�de����[�Y���������Ȉ��Q�����FFvG1Q��Lf̺W�]��!�������"*̖�)�/lC�"�u�f�L#y�=U�뼝�eUG#2��eUo]��G++��ۙS��v�ʍ�\��f���r��*2�J�W�7���Gz9�QT�Us9QV���㕑R��qȈ���һћ"9��D�܎r39Rgb+�W*����C3��-!��%(��k��G�b�wXcL�50B�u��B�;VDd9���{�D$������:�'U9��r2��z;m+c�n:1ZS�(��+��"j$�h�$�R΁�
�5�Ů�ɴl)hNler�R�"b�D9�іZ�̌�39��-�a�1LA�b����\��k�#3�Mٖ�c�frQ֞���׊��&ւQ�������	HQ;������s���ꬷoq���ʨKc9�J�fDB��2�U��Ȩ��1��X�W+�r�Z�wL�Ȯd�u�f��I��_C���D�<I=���C��W�O	�)�Hy/|���tcO|��ik�iW+�h��rLok:ח��f���c+1����Xu�l��zu���d\�_9�"z�����:�c2���Q�qfu�|�ʥ��+�9���os���$*��U����Grμ���~Y��y.b�1��-�j#�zߢ �~S�<��L~r��)K���iy�ũ�������󔎵�1��^���Z�Lȼ�<�|�>L<��j"��i���fT�{��k��[**�sQ�fLr��+��S�܎N��7+2�2�Y]�}ʲ%F+3{;./W���2Vs���/"�{{J�u[��$V��JHBY��c.Å�Q]=܉�b�ݍUyt��Lb��E2o&b!u��j|�SLbc2�R�O��z"�?_[�H��Ȉ����&mk�16ū|놴�u�,�uN�ikj��2��1Jb��Yt���2Ww+Ǝ�����G���5O&4ӾJ��V��)��Z>�I�Y���Fw�1�c��sy,Ɣ�LS���O��N��<��7�ԟꖔ�3KQ�������Y���ז{G�-2�V�c5*���~D �ƚ�⒳L��J��qT�(�B�������I�������Ϗ,����!�K_q�Y�)fC�l|z��Eә#"��7mƉ��#s7R�)������U�KU�oY茍=��sEcr�/2���fb�5���8�\ON�1z�d�LBY,�d���Z>ok<�G�����ܳq����R��-�������Z:��3�y-��9�,��ZT���I���9h�^Y��}�5�5��X�4�$����)�L�ˇ^rʹ�T�KKj�մ�F���TuND����ȆG)}զ�3WiM��/��ۋG���:�宥ĩ�1��b�KdJ��1I�-If*՗��yfڨ�N����7��m���ŚU5�;���?�?=M��j2e=�0�:�~S�Oξ�OߜK���j��-K�#ϼ���o�3��%���-J�\�M1+i+Ýyh�>\<򜓯��;�nEaliL[M4u�l�;�ZR�1J��1*J��Nq!	�0���R�����f���)�m�a��b�����b��yb7�̪��}QY�����m�,�^[� BMy�f�=J����b��.�-�~~z�ҜIכ�o�,�M��X�ڍ+I^�<�|�O�[HA��<��>�g�W�1��dUb�F�����y�3�y-��>�qzJ�ŭYy�����)�{��	
^�Ȍ����R��1+fg_y���7��?<�-t�cO�^����ٵ0�[v�)*[��~z�mţ<��u�9-�%/>�2m��kJ��Ѿ��m�����ּ�m=J���[JƱ����9��J:��7�<�C�8��Zbc5s��:��Ϭμ�ñЉ%$N��S�O���%]�Y���%e+���R�Lb	HR$kx���#�Z��z���Tt�UDdg'DV;+ҹ̇;��d����D9"�ݯ�+K,d�U\�jj��뜞�=����T�\ɝ"��GO#3=��,ŧ+3: �?:��i˧#�i�j�fd��h���<Žu2ҙ}�Μf���WOmUk�Ӎ��5Ś꼓M=䯋i���9�T�GYg�dX�-*��)�&q����s��Q���4����.o%��%�i~r���N��K~t[_>R|\�W�S��%m�~�@��S�M~~Y�G��L�խIŲ5m���4��כ�u�<�����-%�2��'<�<��c
����1jd/)k%*Si��]b3-Kc����iG^}f�n��D��M4�>$P�-�Z��Y��p�s����ȏAOb{_RH{5r�/�feT�9Y͗����oq�3*��G9X؝��b�q��K\�R!)��$0�H������FZ�e�fkzW��|����O<�זi��yȜ�f��Ҧ����N5��K~Q��������ZSXȥ1�%s�9�>I����+�m�}t岚[Zb�m)��">���]�y�?$���y��]qLM*ּ�is�:�imc"3XT{��q3��z�YL��ι�u&�}f�����S���G�g�[���[/:{��]�*4y�zQ�8�:��ןY��x�e���)�Z�,7ז�B">� ����i��u��%�{�-K�\�M1+it�����y\�y��o]�T�f�4�-�yۇ�S�k�:��6۱�Y4�-D��4uʏ$��{V����ʹQH��
����z����᭩ęזi�}V���ZUn�V7���K]�����މyw�3��y��}S�i��y,imF���Y�w�F�|�k�y'^}o�D�?q��ט�M2r��������Ϙ�L�q-���"q\M��0ī�>��<��Ƕ��J�/IRص�!�)�5ŝ}���g~O�%�]35:R�[Jaם��E�N<�C�w��X���8���13'�|�Nq��y\��JR�}��i�߷���vV��1r�����F�>�o�-k�6Ӵ�Z\e���E\�}��"�I��lߟ�d??%��Zbc5s������Y�S�:��6�S�GZZ֚j�WlG_yg��5�J�?���"�>D�w5���U\�̒��Ԫ�W2�+���*�7�s����dr9�����uG!�Ur��jqב4�uV�rn2��{���bjĒtu����8K׵C�;�2��soFr";�ѝUiY*c�b���]�5�T�_8��-���������yh�.�W>"Ui��9ʮf�yz��wk��)�\o�8ң�:��1��{/�jxMp���CKK1��e�KbZ:�|�h�^YԾ�n<W���^4Ś��S�6�����Fu����L��4�[#W����fmM��~\7זmݾ<����&U��Ǝ��(�ϗuO$��Y��]yȕS)qL��#}ye?�?,+/�������:=�6�%*�NRֻ󯣒q��3�y,j=r'&Y��<�:��A2���!E!�����(��1��\8c}�ɭߝC�w%���=�9�+p]z��ˆj�5��<�ܙ�'ݲ��R�J�K头[h��I#kY����x�ò������j��K3LM�hlO:�׌�·<X���q���H>���!�pc��PRF�ѡT��Ѵ����.ֵ����\�ə�F��e�t�$��7v�I�z�;2����ٙ�g9���UT�}7�3��o9I����r""#2ddr��#�Q��\��ٵG4ކVוvF���t�x�s���������Q#��g.g2+�Vdq�����NG��UF�r��sW!��21{��s����̬��g1�Y̎�r�P�9�QV[���؋���G#�2t�ē�g1�y��C�y���)�u ���!7kHML�&� ���;�,f��� Ґ!4�6��1DD1������W*�z+���k
�ӥ�d���&s�H�̍�W;��UVҹ���\��Tr29ʮfg+3��#fUF�c+.q����B(ȁ�D}�w+��G�*�J�x�����"���ޮnZ�g/��-UrE��s��y�̨ޗܨЄ
	�6(��������ٙU�ܓ�*M��3�b��pw��<^�	\�r�M1�N-L]������YԾ�u�ok�xֳ֔JR��My�9��Fu�yQ�m�}+�-��ڵS�F����8�o�y'[��:�宸��U��f4}ח|�h��Y���N�O�a���X���G_���?=Ẏ��*QQVƸ�\*��^+b3�y��>Z<ߖc�<r-�mi/Є4�sT���kFD58�5&�������k���d7��{�z�.�.�iKR�^���<Ȩ!DJC�D*!�y�F���,ֻ���-)S���<�i/�Q����o�m�����L�m1+cMCm�,�^Y�Z��;~�V���[M5Vȵ䟝���\חb��aɔ�*H�wwf_\ތY��8�4������m��X��}�G|�L�f����2FU3��h�\��p�^Z:�l��Z��Jd��}yg4��<��7זn=���zR�Ū���(��-�CRDDao%����s��Vf��ҚSGP"%���;�Fy�g�ߗ}z>�e4��-F����J���S�>w�/�.e㥊☬sO���!ľr���Ӵ�z8�b�J�*�S���̬��/>{��~,�w/�u�,�^Y���qĴ֚N��[4y�?DD�o�5�O�?7�fڪ~~�qjk�^�v�:�q��~�D	o��<���-����J��Z[KJ�֏���f�Y眼Ob|��C��&�.v��[9��ܭ��BU���GeF��sD>��ȓ�\�OU���'9��GVU9][�K�Esd9�Ww���1R�ٰ"�ĻVHU
N�!�d�#���%��պ24�FFS2�ٱ7x�G� #�ʵ��q�����iJ[M%����?6L��-w1��ѡ˖J[�룈�ʻ�]~�����~Y�����V�D������X���ڱ{+3O%�8��u�<��6�ɘ�T��.2��|�6��u�.K�Sn���-%�2��f4u���|�gS�y'^r�72��D������)���͸��y��~ז����%���)�iLSK�C�~z�1��iJr�*6�r�-��F����jإ��9�5�Ѯ��;��i<����ĥ<��Jc1&&)&�F4��z���g�*�2-��J���n�/�&�ꎘ�R�t�\�X�9�KDĆ+ q�|��1[�G9��i�]S2�E[:�|ۖ���<�w�r�M-�K�F���q�.y�G[�߄%�ϟ���iV�Z����?,�;��<��y��i-�񦭑�ij�Z<��8�<��u�,Ǿx奙Mi�is��Y��|���'�h��D#4�����$�.q*N-K�_<��>Y��/%�}�)K����R�������1J-�2%k^���4��<��y��g|�>�KJ[M%�\�������X�NT{���������u�Ӧ:X�V4ӝu���D��1�8'K�Ie���v�:Iqŝ�;�������f��d��	�Z�7e��|�_.�_�F���>S�Z{�'��i6��������M��@����k��ʹ���Kqt�ikj�)P����I���u�,��S�%�-��J�XѾ��[�L�EE�7e�1*[,��!M�z�������>��N��=���SL-le"&1h:-��&u���_��Tm'�yf����v��R�/Ji�4�SP��Z>o�3�y&���;�U�9��[LiM#�=f�)�SD��i��ŦVI�K���������G眿3�쓱�FSM/��h����q�%��<��Ӵ�Gƕ�kQq��FLU1�jK%LR��S"�i�M�8�bؾ7�i�:�K!�)�4�4�ax�0�'P{a��10��ǁ��;����f��ߑ"O>��󏮟��iMbX�Ԯׇ����Mˉ7��N�(�O߭4�-����)�h��8��5Q�y�4ӱ�����bR���u����(�~Y���<<)JQ>��	V�6��R6T\����sz���&�闕�r���fFf���b*9��k�c\���eg&k�U����R�ڢl����(�%lbvTds����I�a�5G�.�x��J7�4ۻ�H��S��%�i����i��Ɩ�4u=��)⒴�2�a,-�d��&ԩJ�+ZإǞw�)�3�,ѧc���J�5�1s��&.)�1*^\�v�^���=f�|�u�.K�Sn���-%���FcF���k��:���y�,�mל�R�*i:k"�o�,�UIל�]yfGv��.�L�Jb�]�K�Q��Y�yh�^Y�Ͼg������bXƚG�z�S�8�%k�TbXB�� �y������0�qǤ��,�U�&�{�\�l���>s�|��̊ު������s.�B������8��[z��	R�c:��D!+zw1��%���Fw�"���ʬ��g4s6X��-)�-�^�~S�N5���~r���u��j�3"��Z�}זi?qH��Yה�[i-�񦭑�ij�Z<���q�k�y'Z��{�%�J�KL^��xu�,͸�k�,�~�{��2�KK�SL:�T�iJt�*2�֔�E���FZ��La�`�}�����Q眳^�T���---k��cLa9iJ���[������i-����fu�{�(�ZY��J�t�����q�}aY���r���̋�+�+�/�Kf�Srg^Y���Z��钕�QJ���=f���:ח��)����K[Q8�f��}yh�o��~�漳M�{�S#�Jjr���������M�kbqx�RT�+���[HKˎ��c>}6��5�?%�|��S#3K~�mY���K�dg$�VG9U�?^~??Z5�3��G^r�;��M�9��iLZ��F���q�F��εQ���ғ�w���LkRe�������[�#�U���u��D�#�ӛ^��+��v硗��8d���F��71
c[R$I�����k�gNcpǣӞ��6[�lM��d��x���v�x�<xp�˅É�d�z^�v�\���"*��U��3���fFG2�z222222"#!���f�]b�I&j�M,�L�Ku�I&�m6�h�39Y̨�U�DdddoFFOd�DDds�####��eted�U��eus#��޺Ȉ��ʏ�|����"####"#-dEUVFFj�DFFGb�*3����*���u��e���ō!��)�ȶ3��OX��s��K�ef��b;+��/�V2t�a��C	(�A!��"R��U���eDG�����H�9�U�e���ܮr�O3s�7*#+#1!U��sٝU�Fgb��;8D�5F�J$:�)ޮֹʮW��Y���#���=$es�U̎Es��L�OFc*5�m'���M�X�-�QT���ڭD�B7G��JS�S�)LC2ƅ�%ג�A.�9���EFG3�^�V�,���GUDdg5�I��"��+�97GL�Y�Xɳ�*��Gn��,ݭ�����&N�h����*9ͻ�3��܎Dg+9�:ٌ�l��#9V""���ڤ�Ȯ-�My��edr*�9�r:ʻ�̥q%�iȎ3�;��,C5���MלE�j���wc��":"'�*�l���"��L���R���X�G�{�2�)���fs*���U���&������4���ZI��rFUWJ}�T{E�<��%���>�}�L�4��DQ�6����4�iW"�KV-��Ə<��O>R3�,�Ϭ�<��8��ƴ��ٍ}Q�b��Ώ��_e갭96uu�ȴҭvťUם�)ĝk�:�����iMcL�KL�%KT��V��8]ܮפu�,�)�N������X�޴Ҹ��kM-M4u�m�k:�G�u��c��yjJ�2�J�ƚ>�ˇϟZ7זgT�Yn:�]i+�im1:����gY���N~��C"*�J�t�eG"��)���39���K�V-��'	B,�	M
�r*5���Fs2�2�H�u{�k���W�"����
"t��1�k�Z�dVDd�gJ��_2u/��;է5Gzz3+�q��_�O~���g�GR�*��F�ZI�,�~(f�S��D���N��	x��u+e1LK�u&��p��Y�v��֖������Ic
e&bغV2�2�37�<��Ϯ}O$�<�Zu�.T�Z�ˊi��DA	|�GRy��5�?%���)�ssL�t�)�0�|�#�>Y�S�:�y��業)�S"�i-#~yf�S�7�u��%���W*_#KSJb����Z;r�[LS"���Q#�}�ިΰ��̌�θm;K�o�,��ߖ���}<��p&\2p^=�g�q��!���lq�s2w;3I�Y�g�[���љ��ZR��y1�dR�IzuÆuYΨ�.��B{*�u��G�M��n�S"Ә��r�.%qk���O�)זu�>��Ko<i�de�U������9Ś��F���{�qr��i�59�9זf��N��O�Q���)K��i�KJV���s�7�u�y0��,�����&�J��)�}זW�|��"-r9Wףe�.WQKU1��*/�>�ɽ��:��ۿ%䪹2�-�W�U�%���*-�b�Qjb�u=򑦾Y���g�~Y���V���f��}yq�1�����>b�i��3335��lK�eRrI������G���?B)��?-�Li�b�J����)�&�}p���Fu���%�D��)s��c��D�=�g_Tq'���^~Y����S#3LƚZ�h�|����{������G9�9*���Q���Rg�-<������9f���-*��b���ƗT���VF1��b��%�����s�o��#>��7�K�v��Kkb�-yO��o�����vM��n�	{����n�LU)y+�<��p���+ G�M?,�Z򛆞y.-���%7��h�"<��J8��5�?%؈�o��?8�W�-֔�bX�d]a�,�m/.Z*U�����c%$LG�L$1M޽��8�w�O%�;�Lʜ��ڛ�_�ې��Qk8ܪ�|u.�G�|��ג�'���O�9�d�򭤭li�~~[� ����$�g��n<���W��֡Ω���:��Q��Y�o<���%j\fkIG\��|��5זJ6D�l�̥�mZ��۷�%!H$�C�Ki;6��R�Y�'��3�����E�t^fJ�:*:9*��F�=<��eG*#��ʮ�Rr�+hȞ�}7Z��]���U;\�B�z�����5{�ԥ.���}�q'�2��-+c1JRԶD���D4�<�KM��Gf1X���F���^[-W�SVB;9b)/z���JԤ��ec�>s���q&u�ӯ9K�-�[�\R�V13k���)JR�)-w�5�q(�~Y����疺��i:JX�Xu�zQ��Y�yh��Y���=��Z�Z���K��}�ѿ<�]Ty-���JJ�b�S^�uO$�>Yו�?B	}��<���Un���*�.?�򜮨�EO~[39ʮT��%-�J��'����g,��,ƛJ�x�V�	��d�)��L�A�7r�B����Y-DM�|ɍ�LC�M�����a-1w���V�$U�HZ��A��
��D��a4�jV]�Yt��UI�8�}S�5זc�q*qr����NkR�u��֎���~S�i���%w��T���i�w�F�|�k�y'[��}�>������cJa�^Y���Q�<�<�ͽ����D�Kb���yO$��-)N��T��Ī,����!�SQ��R�z�}>kkG_yf4��ҷ�b��c4Ң����I�������ϸ��5ן�!����4�����5�e*��4o���Z�����8���<�<��u�|�)Rҹ˺iwˆ���~�KϿ,���7��J�W�[M-m4y�Q�7�g��N���rҺ���Ԧ4�����ޛ�B����\L��`݈0TĢ&(�������o��]S�k�/G+�M1��j���u,|���͕͕�>?�yh�8��*9�yGvڕ���M25v�ם�s�-זu/��᧞qKiMkIM�s��S�8��ڋi334	D���C�-זm�W^N8�-Lb��yrs�,�)ĝy�?"!>s��6�?է4�cJiMK��yl=2�Q6���ZKȤ���*��qt�I�c���!�)Ğy���o��iyVL��qtȨ�$���r�3>{��~)�j���^Y�S�j4���.���ť�C��h�8��o�:��6m�7Ƶ�M4�E�<�ۋ?K^~Y��Ge��?i������-����O�\<��?>�L�BRw'p�1�Ht=t)�����m��ّ�b�sT"��1������}}F2�r&�Y63"���#ٓԮr����$��JA'ii�%�(�t�G6g-m3�}S�����\S�(����Ԝ=R#1��;FeEFs�ʗ1��G�����V-m&�j),?;�g���^�Z��E�LFK"Iآk�a�T6�1�=�?�f��}yfG�|��74�'II��V�J"`�{Lc%1D�>��ߓ�<��眳mm~z'S���e%m4���4��(��.��4��].��iK[JiZ9ז�5�μ����6�~Z���Z�IZ�u�K�g^Y� G���m�T��5�V�j�}����[��"�]��eh�dgoX�z��J�.�Ǟ�ϟ-k�1��v���M-R�\-L�	L�1��.��n�ks���.�Z�c���Թ��8��c&��Nz^��uQ�K���S��G�M�n^���e�<g�gl�����Z�ޝ9�:+e�&�0gn܌5X�`ʲ�*̆,�gI�ı�1�Y��d�����zR�v�c6]�^��V�Yd$kIա�0F�le����də�̱��ǋ=.�t�cfVLv������s��n����a��gE�-�v1���FZ��w��339ə�Fs"�*��{39�c6�r�339���r'����ff2�ݻ{mL�k��r_3�����9$����s��==�1���v!���#���ee�9N��eޮW+��ȮdVVr�#�ug;�̨�s��U�9���29r��=}��Јە�U���R=��ŝ����?�%<('���!����	H��+���a1%q�����	u���Dr�;�"3��T�7�Վ53��hs;Kr���uE�9qU�͵������Ds&��JsR/F��J��b9�2"��U|��s7�+�]��m�_bT��~�'�+��5<���_)v�Ϯ�:�]І)LS	��B��g<�g+)�k����ќ�җ����,��\M � ��$!IK�!2%0���">�uFͥ��1+M�+,[�c22�jO����kG�r�Ծ�w=I]�4�%�+cGR�i�ˆ����YＧ֗���)li�ϼ�TnN��זiݥ�z��1Qli+�<�|�m|��o�:ߖcNϢ�⵬J���%h����:�����R�T���ZQ7S��ԯL&V�{�Σm�g�~\6�o-/1���-��s�&1�^Rmx��J�e4}疍6������)�JT��r�G\�Ԃc\S�y�7ז����[��ĩ�tҙm4��y�ˈ���k�u��cn�.JSY���kiZh��,�-o�?DD	ߔ���)~��b�cLV4ūG<��y�J���}r,Oq������\�M�.T�G_y��qo�;�ԯG.��27s��έ=R���q��h���8����yg[��CN��Қ֒�c1�}�<��>�}yh�^[�	~p����J[V����#��Y�)Ŀ�"~�&*��%8��eÓ'	�'T ���p�Z����<ZsKf4����<�|�ˆ���y��c;�&&��Ɣ��N}�יt�3{�8⫝�%�o��K1j�N27�����T�[�=�~9=oʷ�>̞E�I�ֶb���P�]�5ŝo�G[�͛y����֔�iL]���ٷ�O5�חh�ʗc2qqu���yO$�n\<��GZ��iלR�k�U���:�mO�y��Oww���!���1d�n�W�UʌΨ��z*��Hh�S�rl�Lb��Bv������⺱��vt��s	���g���{�D�	�6���SY�҉���/R�s;�|�Du/'Us�(��=�B�!�Y�;�* ��ᑾ%󉺦ij�UIi������_�'�X��М�ve��Vb��U�Qk]��8kjq'�}g�>_�9<�kT����%t�/&�8�Z��b��i}�K(�~\5�<��{˥ڜ�)kiM+G^zѦ�Y�yqo�:��)uk⭥�ib�^v���,�����~S�X�iS�Ɣ�eZU����)�&�rμ�<��=���8Z��M\e�:�z=�%-)u��Z���sE��b-w���s~y�>}�ï��n��)K���մ�9�6��duoETVTD��z�C�nJA�7L<X�]�ƴ���. ��]������w�їѓ�s#[<�t��T����os�qKf-J�1���m�ᾩ��"~~v�ܗ�-.����-��7��fi��u��o�y-;}>ZV�1Qlit�<���uO$�^Y��>�[�ֱIR��Q瞳���g�Y� F�.?%��<��1��J��M���~��'_���ԶR�L�����*mQ]�Y�Deeq�;�����,ǼqN2R�i��gϛ3�����H�ݯ4}ח��h��Yה�ߟy�S2�[�F��Q�#H!��b�5壭�f=���J�5iZ��i��yg��~ %�?.������.��b��+?)�3�,�*<��9gv�]񔔱q��i}埢�~�k��db�7&ZHn
&�	B��	���>�6��<�?%�y��M[M&��ť҉��#���q�����h�����}&u�h�G�Ɣ�4�^��u��|Z:ח��)���x�-:R�iMr�I�>ZK�ebL+vNR���~t�<ݞi���fT��4���pߞY�Tm'^rξ���ߖ�%u��T��5��(���&nb�Yv���s�4�����$w�1����O��k��6m�ފ�SZ�b/��|W3WF-�^̊�G�z�8���<���5�?&4���N���X�֩�?;�h�_,�c~Q���Zy��Z�2��.�G�yg���G�rμ������f�i]i-)����~dF�v�ϩ������;�3*D��K+2*/��1�j��ffdF�Ug{������6܎dE#����"���k�_#a�R"Z%/n0�lGTĤ���\h%3{t�J%dKȥ&� Mb!D����X�-$��[[���D>|��,㯗�NObZ���K�s�;Ioϕ��}"##��V)lbT��1LS8�\Fi��N��6��].�Ɣ��B�	�I��6��4�Z�dS���=&��fy�qy�1��Z��ůKk�����&>�G[�η�m-�x�V�M�UZ����F8�yO�μ�N��N�.�.Z���Y��'Z�Φ7�6���]�4��Sli��yh������J���)k�;�\�1�:;*/����q?|�y�,���r+��cM>�c��?]d4r3l�e*�g7�/������9�̌���������\a�%2�)ju���w��n3"z���ϾC���%�L<G�JW��bT�'�~yfq��u�,��y,v6�|S4Ңض�mLs�6�u�-y�����kqVִ��W���9gS�3�,�<�i��Z^cKV�j��Z<�<��|��ߔ����)�JT�1k�\����ս9M��J�i\K-�&�6e&7c�|�|�q���Ϭ�~}�%L����)�6��ƢX����Qk�D��6}�Dcm����k�1ݼ�&%��խlV�G\���LDE8�>IןY���;�q*\]r)�4֒�����7�gT�a眳�|��n2Ӥ�L����^Y�w�#������h��)ƔƧҧ���^I�&?F�ԉ��F�7��/��KKjc�\ᦟZ3�,�ʟ�K�)t�Wx^��ZU��br�ldR���u��t�L��:��F��i�⪭��ض���)�6�N��y�6�i�ʊU�1*c�o�,�)�ƃĒ�Q��+����5��1�����d�����q������� s��<�R�h<!P#�'NDRI���Ag*��ܧW�g(3�r/t��v��:GwR�5f�S͏�E�����������r�v&��O˧i�3�q���ۧ��c,b��c<3��1�S.��=%�\<�d�L��p��,g#�3�,a������-���L�.��dÆqd����+�<����f��a���X�1�\lp�.����3���ώ�/ƶe�GYӆLe�&ZD�TI�%�ҕ��1�a[Us���fW"+2r�4�UY�F!�$�M4���k�m�i���L�4�Id��&�Ha�!JA�W2%VEFFG9r�3���#""&s*3U_K79��.�-�UFFFFFFDDddddDD*"��QQ��2�###)N_m�4�4�3v��J��eU9K�r���dE��.���&�^r�7gr[�̇wd�T^����cG�;�eD�[�9Q�X�Vf&"�""��"��r+�Y��ʨK��EEX�u����f��r+3%fjʈ���fr���+#9�Ue�T������srDfsFj�FGfEG.sH��U�q�2��*d�Dg'�]�TDG)̾�r�:�W���1Lƨ#�Jc�Jؕ�DTk��y��*3�1D۶R��$)J����%��B�ťr͵l�R�L%�9Un�Vw3������YX��3n!s���c��W�B�kK��g��n�#+{z��\��v�G39̌�;&��U�d�s2�"��,��ݭW3�F��W+9����T*6wtr*!�n��!DY(��A�b+Т�B��ib���Y)*���eUw"2�-���fDs��39Ȫ̈�Ȯs���f*�/���FW#�}�ː�ّ�z��]]d�/.���>���ЄGH;)����r��/��U�>!j�v��.�5M�����䮲�e-����'�R>s�:�<��>�f�}�˴��j��.�y����h�#���\��JFm*��4J��e)V���x�����Lcg^U�ƚV�K��./3*J֖��Į�����h;Y��/���,�<�V-jҩ��.�:�|�|�y�,��}-Gco8��i6�֒Қ7�<�i�y�����4۫�K+�-KZKL[Kî�f���:��?@�$�"V�mґ=��m���fW+3$�_fs3�\ި�;���Z6�Q9Ȯw;3L�����g"2!��W+"�W"ѱ�SrCX[%�7X$,����*,���w��U+72�w�Ub'+�z��ދȬ��W9\���u�^x�{�B-�s�O���.nԖ4��,h�������~�*�.LS��z�k��q��	So��g�0��Y����V�-��w��|��\dX�eEh�]6������_I�ߖu�y-�ڒ�Ɣ�έT�V�9^J4�y/>�]yfݍ�8R�i���u��ϖ���:�%����q*J�K�N4����Li�<�y(�^Y�ǔ�W&r1��m)�y喧}KH��!;X@J����������F1,ߟ:�cm���Y�F�O�f��ȈAMmQt��1Kdr�/9�F^��9y}�yS�=U׌����Jd_BC&� ��6)�&�^��v�*�9u^����w�f_d�q+�S�1�L[���.I�nY֩���?>�O}�R�YlԩZV�Kb<��ͥ�(מY�yp�M���Ɩ�2�ue���L��O��N��w��%,Z�J��#�9f>��O5�Kϩ�����Z��f1M4h�^\E�yL�b�Y34Dd��ns��$��RR�)����x|�>I�yfG�o�;�����~"�I�|�e\�[����מ�O��u��D#7Q�/���)k��4�bZZXy/��(�F�Vf�\G^r�m��b�l��4�ka�����/�� �������0��q�1��i3�h����M��Υ��k�,�|����J�Y��j#�=g�Ǯ�TxP��.)X$l����ӋZ��:�_8���_K[z_��'Jϑ�MU㖿ҙ��]h�b�Jcg��m4埚����yf�m?yQJ�Ƙ��Z��Y�|����ξ�����i��Ym2��KKGS�'Ϝ�}:�y�y�5<�T��2)lU���,��֏7�ЄDk�~Lh���K�1l�������O,ɩ�S�xR�ݓ"Q����Fَ���1������u�,�:yī~sSzH|JeE�We���Vb�u�,�����^Y�Y��m�T�-Qu�����O&|�}O$μ�M��T���1J[�����m�G^n�5Q䵦��]ZRƔ��M%��;h��gT�c�����"z�)����ԤE^fw5B+���;��w7����Z�4rTV�=ȏoH�g�����EU(�R�J��RD�A�	�:��yى�l^�1;�����H�wHY�YY��
ʮz�T�̍s�C���yvm�|Z��ůKk������֖��S0��R�+��뙕}������;ȍ9Şy�1��u�JS-T�݄��������lHM<ǹI����>�u�,۱��
k�S'Q�^v͹N$μ��>�i��=�f4Ʊ,N��眴i��<�G�u�,��^r'�9���f�����,�uI���y�~K��&|S4�&1M)��v�<���U��֯�����Y}��]]�*/�uÏ�Z:��4��*S��k=�|�TWt��̙����p���#+2�="*�ef��tUn���cy'"��u9-F�s$ī�,��396����"B���w�BؼM�8��ڍ)���,�nZ<ߖu��%����Z���ձ+��<�f�Y��a��Y�|qN2R�i��9tï;f�W���Kϩ����e�-���F���9q�'9g���g��dz6�Uښi�iY��Qs붙)T�"�1h�0�/R�dx���S�{�}$��Y���:��q+^+-�2�k|��C.��ʬL�dUs���������Լ��>��>y�V-��)i�������DDD[�*2N��j�KGcϔ�JcS�g1��甍��Υ��u�,�gͥ���R�ֵ,��������-��~TnZ���"Uli�ңM%�ϩ䟡�ڧ�Ke-v˓=͑��R�5����ȸ���8���y��6�o�ɊU�4�y�|DKɂQ���ܔ�&����6��<��:�kn���t���KcKSG^TrM�Şk�G�}fCO<��%�ȕ�V�u��q/o|w_J��23%��0�HCp@ȁA�3ˆ���4q�K�)�ebS��מ�f�Yו��%�?,����uLR�r���H����m>it[JslR�X�eT3�+3*~?^�T|�u/>��ѷ����LTƱ6��X$1i��1�#	{�_^Z>m�:�5�۫�dӑ�[M)li�I�<�mmh�Ϭ�c~Szm��ͥ�-���b�:����8�g^Z<��1��Z��ű�b�,^}�iQ�:ߖr �%$�>�xzwp��2���Ž����;��Z�nɆ+3g5L�tv��t��l����Y��qӧ~g
����M�i�ݕ������4�Vb����,�D��Kۨ�����1�u(�z''�9̨����"�zW:�UD����Fv����FP���Ja�Ä�P�^����j^L�I0����S,̺����K��%s�U+R�Ls�<�ڒ�G�JQ\�+oE�<��f�rfq���ᴴ�o�6�l�µ8�J����^�Ȇ*4qJk�[����|��yg^TnX�~���i�bX�)�ϼ��8��?&>���~[��%��"T�OY�ض�֏;�p�>Z??>��9fvR���LS4�i*SL?Bs�":��?7�ga��|���T�)�j4�h���:�1�認�I�ZJ���E,�&ik���Z��=�f�\�/�i�����O�J�(��R
�����_��(\�Ts*(m*�Њ�搥���/�J�������J�o��z�����������������������O����YR`�b�U5J�Dd�Z4�5,4�ɣ-��4a�4hɆ�MMi0�h�dba��E��J�h�1&��Ѫ�Fhb��h�%�Q0�ZFMKKF��F���Ѫ4hXj���Z4�ɉX0-Uh�+F�0iMCF���a�ɔdd0ʰ���a�ђ44�F%diI�)i*��#F��I0�#$Z4CI2���E44Jщ-)a�F�IXb�E��C
dj��	��j4�5�DѩV�BhjI�Q-Jde#"��-J�ʌ�$�*hb��)�JhԲ5V+#��djF�%����24�`�&�D�0FF���YZYFSI24��j�����`f�d6��E��f�U`eFE�052i
mUUC������(�����bP�?�����P>���J�% ����{���@?������������?�ο��BP��~��o��������O]	@:y��G�����J����z������1AY&SY\ݽ�ga߀pY��?gݐ?���a�>�Z+��P ���W^��ج`ҵ�Vv5�v�             �N�l�E�
4h  ( P T< ���D4���S]�n��V��t�ݭ���s��u�v������R�(�y�;eUW��GU
��=�@;m7c:�w���ԠV������t��(G�D[�HT�X��;�`:iʇ@����S��C��z� O{��ֽ8�����D�[�9v�Wi@�U�U�`@^���먴e݀]���V7`��ϕP�w���|x� ������t�:�:Ū�Z�c����  
�n��y�h�uuc���t�@��t�Vޝ򶂾' �{���A�=�6�<m��O|����xf��nXj�=罾�())\���:�G��즪�ϭ�z�qC\�]�ԩ]���hU��t�h�@4&Z�V0��C��cg� H���ק�:��;������vt�:M=>��;@> =      �5Sٓ*�M      %1f�*Eh�4Ѧ& !� �2�I�E       	OB�
��&d`&& ��M
4h Sj)�OS5L��(%R      �}9�������������N<�����
�훧�}�PT�$>aAS��#��~GZ�����?������?��b�f�����MƟ���r��
�r�Զ";k��~�};��ݾ������L�oy�^����WF����B�u��e�Z���u?�򓰷"�桫����������ϟ)k���D%]q��|��>�ՕBT�^v�7j�vɶ�U�:�j�,��{ӁN�/��$�8����]*n�]�����:��e���P���i1S#B���!��[�������K*��W]-+�^T�e��\�b��Ykﾗ��x�+�1���0e4w�ݿ��{Ŗ;qp��|K⦄a/(S!h��	��^�Rg�*�	L;g�Im����\ϩKA�x�]��Kw���	9I�^�2��O����I����?����O}��)˫Xr��KQ�z|��T�������g���ØB혋|8�}ʦ6	���O��.�l�&ɲx��6Nd�"�Z�de��ugZ�vf�u^J�;��TƋ$���1�i�]�v����;t׏:b��3+�M��b,�I�0��T�Ԋ)S�M&�T�T��m�n���q6��Z15Rl�Z"ѷΤ��6c�N�+�jF�뉲�#i<e9�����[�=mZS��k�ޜ;9N#��&&�np�+CI�`��}�cʔвJV���Jbk����~8vp�z��n�l�ƫm;m�����4��uC���4�:V8w��i�-C00禑�om��������1jJ��i�C�е1'T1l���n��0ɛ)ߜє�2��R�,z�)N��&�2��*Ty�x�셤ZE�ZM0���񳴯+�lq���T�u��1ZU�4�Ҷ�벓g��d�LLZ�h�xڱ�0�8z�U�[N*�Z;�4md��#�ۧm�WO�+�UXWn�=ᆛq�G%1�Lr�m1�'EM$�L*�Ѥn<�43Z4��F�#RqҚ��NN+pp�8�h�kF��4Q�kI��w�4㲦&�6���J���jN���4���F�ચ�:EMh�64��I�٪��LM&���T�*�v�cM�Nl��a���F'y�i���84k+N��js�D�N��w�����:�\XP��R�Ç>�y@_~S��;ϑ�p-S	QYCT	���vd�.���4���w��;��=�ş��^���x�Nu�ǅ@ֻ�=ӥ2 Ĩ�A�L��&oaZ_��Ϯ|�y�2
tyo��22�yv"�i$�x�B����W��|�X��EV�WB��])���34:>CILQ���fV,Vd-f�圸�:[�;+����"�����LT_B/]��C�X�B�g�>���'���..`�,�}�؎+YN�S�fC��;�3��qS���	�V��O52��*���G,N��t[��v�a~��Y�%�NK�|Y9Y��+�]�,����y�K�����\���E1�!�TQB�G���d������
D #Q�������b�C�,�y|���YW\���}D��A�4Pګ0�Uaqt>���L�TT��+(��Q1{� C�yG�p��x$N�NA )��D��
	!ۈ�3���W��F���;R�ۤ���������M��ز�0d��z�1���J�%I���ȉX|CZ(B(\�7ܳd��b��\y���|+�%t�%@� ���9feIPA'Q׻�^M�E%-�����}ˮ/��D�U�h(j�X�EU���΅�!H�v܏�2�'�9��.��|΂s2`��D����T��Β"�(�s��Ai�Bb��K
{w���!���_
W�[����T��!���I�1�=��e�8{<<̧2�|�{�I]_�,�s��"��}8�;�G4l�S��L�S�F��\v(\�RBp|��Y𥜟*I�����^V�B.}>��o��T��|%M��+,�!���'�c��pS>�S�T�V�E4���>�R*��_|GR�x�ﮐD2Ҩ�Y<�amR�XڙqF��q��.q�rg�����>p�AҦ�"��P"g0�>�<؎�s�39��ν��-��-�h���1�cN���$��3��<�X��*2Τ��SZ���wF]6��d��U")�qs+�㋊e+U+�����B��,�d�YS��K2�f&������t�)���$a�x����'N�����qP�!��kw|!h�:!+���y�����*�W���}��<�^+*#��qQ���4P�/;��"�|xa��T�x2L���5C���u?���}cM����w�_������"���o6�N\�W�l�S���B_Ly߉�n�V����\d���哉��-gW�CA�TSH�tB��T[����8�G�ƦܮI�pJ�abU��]�������#�I��/B�\w��?>j^��c��r�|�;��t��q>��I�N�ab�Yӳ����5j�9b��,��YyÒ�Wd�&,uduaj5b�ďG�0�ֈ"{H9%eH<��5� �p�<b�Z�Qj-E���L�o�=�)8{՜�A*G�}��"|B5Ϊ=��G�T["�n�VFZ�:��wݾ��L�
�#(D�����}����3(G§*Su��dD* �6%1�gzEG��^]����̑U�r�V	FK8*�)��������`i�};��Fu���AK˘� s��3;�p������w�N>��/ڔ~N�� ������C$uK;$����ó�}_*�',�|w�﹅��DC��* u ��L|}>�]%H�$��.Z�o}b���fqf!��CG�V|�Ht�˴��f+��:N�n��s�&���������D%C.�Q+�`5L!��I�|��Z�I:���w��}�x��B
n�����0A��D���YxK8�yTNUFXZ�YÖNq��sw;��.�$a�*E:1�:�.?�k1�����:�"Пh�0����]�9J���,��F�L�<y�B^�2{��}
�"M���o{6ˊ\/� ]���{^��cX	kFj�<2��>|u��'��TZ(K�^8^�N2p�5��>{�	O}��^HQ��RUB&w�~�*'^)�����1Bˤ�8.�9������B��`a���%|��-NyC�BF�)A���@�ǋ%��r���.̗u�_"ub���`J�Ѱ��)}�M`�"�f*��V2�`���A��5�����������h��,��*���+��a���?������a���������~�w��F��o��i9y��wwc��^�x��'=ۑ�Ktǆjܸt�%7������!�M�ǟ��s�h��Ͻ����h�f�~>䞥J�GO?o=����|�׸��Ie��t�]/�&�y<����ɒI�]z����.�Z�.�N;��K�M.�K���K���K���t�].�K��N�Le��t�%��]��d.�K���t�].�K���PE��G D�1APC�1APC�1APC�1APC�1A���(!�b���(!�!�`�!�7u �b���(!�*`�
(�� !� ��("b���(!�c��#�1APC��ޜ�!p�y�)η�Θ���t�C���S�ҝ[K��u��N��1�u?w$UI�ivAm2Ie�_U��]8�:]2U	t�S�Rҽ�ĺY�:�.�)t�y�)�_�u:])մ�K��)�<��/Ժ�.���]%��͞t�]:�t�|�t��
Py���ߙ��)$�Y����/t���-�)t�y�)�\�i�uT���0�KZv��L����b�K��R��q~����N���]N�L��K�Ӯ�J�ΗK�
].�p�S������}VR�t�얊d��`���t�K�ڦK�;��ӳ:Φ�,�],R���-�K���t�].�K���t�].�K��-�I-�B�t�S8�K���t�].�N��*�K���t�Zl�f6˩:�.�Œ�d�[U�8�S��]N��E"���i�����t��������b�m2ivK�̅����t�C���j�T�B.�N��*���ܓ��rG��].�K���t�].�wq�.�*�].�K���t�].�K���t�].�K���u�m��t�].�K���t�].�K�:].�K���t�]��d��d.�K���[�)��Y4�].�K���t���oYl�].�K���t�].�K���t�\�J�B��$��!t�].�K���t�C���t�]-�}v K����%��,>�t����n����绩;ꢼ9��ϵocYTƷS���f7�͓�3��.����M���P�m�	퓤Ik�]�ooT����cd��v��I���t�].�K���t�].�m2Im2K��������o����wJ>9�<��v�r������95<���^��wf*7�[Z�t��&�'6j���gz�����}�+�����	ғY��λ����M��I*^��f7Ç����Poq�`̯��u��F�2��eI�NN��a��S�ؗ=���r^~�ա^3��~�]����n�o��0fĔ/�v�w}��ӡ��6<u#ڼ|;�����x3��%^w_e���gñ��%%w����)g�9�s����_Dߠ�|<�oyZ��x�~��w޵b����gT��wr����U��&��^�ڍ'Oy�վǻ��>j����'/?.|���K}�N�ݹ��:�[ӸNg�s�Jyd/���z��gn�f{�|�G�Ȏ�=�
+���y�O�U�-���<����wv��C)���5�8��o��s�X[�%��t%������m��
�_wwr���s+wv�z�Dkd}�;W�z�K��Y������o����q�N���~J�|I�`�.f�v锺]/�uSO�fMg�{�ȡ]��+�uܘ��N��Ԡ�0�x�宕���NK:�s���M���-��><�O�.��i�f)-�괗�;�T��<�<�ܾuy�{�o�#�{y)3���r�rxv�f3�[���~��в'��އ�p������pa�hù��7Ǧ���	���Ф}��\�ēZ��١�����,!�f�T̰��!�1f%�|m�3s��A���ktwD�xx���0?G���s�^�P�].�K�2����6���|��1=����㽯�Z坒I%�C})/���:�����zwwN�{�:E�lW���]��w2	,�e�6fI�����w�SU[�N�غ��"��앵������3�wvi�����\��M4����>�7`}����7Ѝe�>1.����{�5Ԛ��5����R�o���4�<ʝ��'z{�����Xp��.�%e쫺���}0��C3Ԡd��,;5���E4�����c��=��s���Dڄ��q`�,'rGǙ�F��F-~8�
#�9�1�/"��1.#�,�|�������S��%�{{Ʊ�����4��^�x�ǀv�"�-!/��A	ܗS��{����w!sKt���F��p�2=�!	%�=�������������-^� �@�7{�om�ۓ��̛�Gf��2��I>��h�Y������9�� �>����gN� �����o�7���r\��n6I��7��ݡ2zX�M���8p�AAx�8�rH�P�N(��6{WM�6�i#�_��"�I-z<��s����|h�#��Z���o=r{����P��B�a��8#�> уG�c;���%�<loy�)v�{��vb~2n��0�_�;i����!b0�㥞:Y��Ϗ���8h(�JQw������#�����]�ۢ»�?>0�O%˼8PA(ЂA �<b������Y����Eo�\8�5�חwit�wy��u�����C>��� ��=[ڮ����8|j���b76��X�]�+��u�y�n���Ҹ���ӳ���B�#�OÇp�0���m���$��!���׽�R�Ӹ�gt�wm唫;ޗ]D�� A���N��ώ8t��||1�<Y��ُ^<z�׌q�Zv���ݼl�n�].�Nɉ#�cU~,��QI/y/H�K6�'w�7ޭ��l|Bt�>�Ő��Y�ӥ���Ni�Ru�µ�C���B�z����ベ�I'ޖ�����!tGH||||||Y���aӧx�!C|||x�����3�1g>|�,t��7�33!m��=�f���?Sͅ<��Y{���xs���o��g5����.K��M�{�s��IR�j��3t�x��B�,���t@DA�A`���Dٗ���S3%䖺{�w���$�t���˥��t��F�g�S!t�qOz���Kz����K򭓜k5�K$=��^��i�>7��~ՙ��I�.��C!t�].�K���t�Im��p� �|A�x���i�g��<p�N�C�N�����d[����ϛ��nv�r~��g�p�T�뺖#���] �K��:����N�a�K�K���t,vae���$
8p��!ᣤ8|3�0����Çp�t�� ����� �6n�n��Y��fY�I.�]�OSA%�{̜�5�tԱSY���{/�U2�L��-�L�S�����v�@B0G8@B,b:X�3��t��ьd!Ӈ!F
�/wr�����I-��/���N�g]Pɻ1M/ܬ=��Ν�X�n�< �� �� #@(-�ڸ��mv۷m�6�ێ8��a��(!�b��C8Aowq<:S$���Mf�wvI-�I-�.3��
�)�%��D��T���:t����ǎ������Hx�������	%�����be��t�{���
d0�龎��w,D���8xA��y�~??���Ѽm��&����m�-���<�8xpc�g�н��|����]�].�������J����E��;sV|C���F�R�v]/�(k.sTζI�8�<5��8�0.�{�&��L��ٜfql��<1�xk�W{U�y���>�܁}Ty��/��x3�7G{�|<?x|3�ū�vvi@��tl�oww�f=����=�Â��-{��u�7Z����'6t�}��7ޜ ��K+�toR��"�<�޵��S%�${�.��ޓG8��0p�� "���xPF��z��Y{��.�e������S>���������m'0b��4GA��8b"�Ϻ&�t������K���ݾ<�<4��̹��N���^-�N�wyèAa�4�|3���!�"��cg��ϯ�ܸ�q��oZ��� �Ts2R�{�;��8�oSΧ�P�]/3)`�`"���(!�b�(��wF� �� "��RXW�����6z���t�]8�j���vL��ʜ8x`�q&ը�W���w}��e��H�]�Χj�w��ۊDN� �[j�M���Wwv��Kqm���s����8v�ҽ|wffgo��,�&wC��,��љ�uY��@A0�APDDV)��J�K���網rʗq��'Q���/�r���^��s��{��$�a� ��ۅ�I$ղa{�I�����8Q�A�C����N����\��֤hჯ������������Ç�~5�Wwv�)=��7��ɘ��I��yvq��N!�ú;��u@A`B3V��w�b<t���{i/��g�莝<xCM�Ѳ�uH���F�Ǚ�Bd��0���Ȇ ��ui�+���x���5sƏA���t�].�d���l�s�d�7�q$�m���)�4�];�!��|���7/f{y�q����斛+c�{��~��.�$+�H��L�ӊN�vݶM~-"�e�].�X�C`#�=�ә�\.�m2Im2��y<o��w]$��"�B��B���%��$��������_�H���Ǹ��/ww_g��p`a�8@ƍխ�����M�{;�6�{�F�Ի�C���������1���3��]�v���!��׈��������?��"k7�<.�|t!`�(z�e��{�z���4`# �@C��yԩs�fdP�n����8=[���h�M��̲�<8p����1APC�t�K:C�!Æ,å�><1�1APC�1G4hA����x�gǋ><Y���B��g��(#F���(!�`�8p�APD�1APC�1AQQA �!EQ�� �ÇA
�G�>�}����J
�S���*��R����q�>�Тt��*�y=T�/����Ox��.����`�䃤��X��X�Y��f���BN��e��R�%M%](��F��xa5���1��`ֳU����ci�d�V�x:�xAԞh�\�ȯ�P�U�#ҩ�Ğe^`tN<B�)�
�T�RyU�S�]�w�qWd�
u�|LSbz�(N��ߍ�ܓYs��q�ʑ�K�MH��U�؄��G��M���b0��h�V�5f��&�c��Me2��:��0�]jWz\Uz)�54&�Q��`֘��OGh�+���K��H;�xN�h�]��)���%�%��ST�̠�<Ԏ�h�1Q��	���*�S4���׸t�Ͽ����I�M�d�6M�jmZUI�ۍӶ��ӕ0�`
���c�i��b.ٵ]��k���U�]Pm �32څ�[Um�̭���[L晵��D���,�A�Y��Iqd$[����*Ve�kv�Rv�V%f��m�\��3D�ڥ�Bǲ:�;a)	�%lؚ%�c�EqR
#�qK3��l�"���i���Q��<)M&��d��6-�aF�Y��n@N��Y`�\X�, �Kk]6�d�*�72�H\�#P�)A�f4�b�:-�Hٖ-h�AM�m6�R��b	�~;���j�eq{+�x{��������_��V�ˬ������.\##4�+
%"�SU�h�U��c�f��2���ø���y9�-N�m�s����z���Y��/���i[Wq��C��wCˈ���Z�7y.,�������_���v��D�/��.�^�	^������̇A��|G���ѓ���	�c(��5�WN�{����=�{���R�m�&mcG��Cm�+u��_i燺wұya��'�^"`�İ�:yU]UQ��<�WsҼx�֙ Ӳ[�#������M���+��Rf~K����-����Y�C����7,���U����Fԥ�����%͖b�.^���Q�����;Ƚ�d��vD���uv]�d.]�ߏ@��eb�;�`�ޥd��u�}��w���g��w�]�j��XC+�u��ª�P>��,�f3�֣Q�]B��UUT��������<g��̌DY�p�<�6z��+���R/iY��Rw���^�J��*S���p妓M�m!r�r���W#��\<��:�_����G� ��0_X�k��>�ӎ�]{���rV�T�񲸵KXn���o0s]5��}q�\���Gr�M&�<�R�X 1UT7ks�8ܪɆR0��c6ˇb����"ZMd�aH�Rj�їK��Y�u�h˓ �V2������,�!D�%K)�L��1������׵�K��C��>}/���H7��E�բU�v�hm�;�_}�Y��_��y��y��o�$���Lg&�w��z����]�ҽ���}WV�R�w�C��q�į|�Գ�����Ř����]���y�}�b����ƩZ�Yp�C�a��,]�9���b�s�ˆW���
�"�v���<%�6J����X}���>*�C<�����:��	�n���.��$չv��e�r�*�	[�@��cY��R�ni�X���]�i�;���޸�xHb��2YNA��WlPn���#�̨}��~�����$"�Ũp����Z����V��*9R\��w�%gw�������n�j$-�`	���oH{��[%K%��!���,@�� ���00�c��֠��>��^?$�y��g��,w��v(��*��$����wK������3A핺��tt�IK��}/��'"��'wS
��W0T�Z���#:EJ ��=�Y��s����1�uxC+�u��:�gxz�z�7,�9�ӿ�]�;߭�_w�]�0�	$s������LW]!�a�B�-���I����Z�;~�����H����6���1�K�;=a�����@�.��_8K��a#?x������,���q�>��B����>h�0�}g��:��{��,���a��\ω^\D�Z��S�He��Xw� �%��|�t��Q�UM�.16�j)����O/7��O�#���s��Ě�[dV�����a��C�?-*�n�������i�ڳ7af}��+����Z����'���^���&��uoB�]D݇՘���&�Wf�E6�:*�u0�ТC�c�`.���]��V�MI˙�;Il��c	t!Pg%mc�]��4c6�6��Z�UY+]q���5.
�c,��U���w��z�噎�ٕ��w��.�.HA4�A�t�"��1��R۳���8���{�Od=��ĢI�n)2 �l�q�}�_��W��W��Գ������,���]���/#��b��>Q�Э9`����݀K�*|w�{�,@��
�[�Y�!g���UK�����v��iV���>@�u�6�������.ۺ�g���W��{���{���<���fޤ
�ip�J���m��߽��xiH$.��!u�^�l4`D�g4��kVKvtMq/I�����[�-�[�|7�5}�V�������\�%Ir�U�x���q|����~���v[�"$-�����/v��iSNBE����oIX�K^���e���|>?~��~�d��trmm�RК-*�nZLg~;���;�J���~�!,Xcn%����u,l����?m�"|+���I[�`_��~%UT.}�puߏC��Sr˻jK��M�;ߪ_w�]tf!%�u#}\�����B�g}J6�9#�=�0a!�Whb.�ZN���M�ܯ}�g܇p~Fy;��	���b��
��
�vL�.�9�w�]�IY�x��r8]2�g}+�?�w���3j���탒�r3L�t�_a�T�5W�嵅���+
�g2!������G��ӣ:��k���z6�X��L����Z-�J�eb-i%F�f�qXq:FSF�I1F6�hTѢ*a��bh�L%4hT��0���L
%)Ի�����p�: ���ҵ\Z�Ŋ�*ڔ��I�n+�\��Srmj��.KK�,ĬX2K1�/:Ns�L�e�ʥ�h*�@����\&��7%���;�1��F1w&�!��#�=×�c�D|���wB������<�����*��2�ԝ,LN�4�������		9���"��<0���_<�Uhi�I@���ȝOG�����,T]M�`�8��9�i$�Bt!�b�!�{	�I���дL�Fm���K��˜暫u�s���v�9�r���0L�M��\� ts�� Ύ�f]Cs��sa��rSX�][f%�\m$�M�$ �r֭ct*M[q���3c���Z+[+lB�X�Q�mj�)� 5Ҽ�SF���[f��s���홣)�[v5�劊imԦ�eBQz���]�S@4����9�I�g�iM�,����BKlk�,��V\�1,e�*�`V�X�q
�s�,�r<K�
����4Кq�3@���Yf�K�nV�a6��J��*�9��!��
&�K��
B	B]��!LQUYtC	F6#u#���e�Frl[�۰�r@l�^�]p��GF☄c�mi��jV��G�"Jy�'$g�-�iDJ�f̳S`�U!c��B�,-tx!�H��M(��4;9&�k�f�%�v7lk��1�b ��JCM6�b���HB���	5Uғ�S�Rw=��)�T�N�#�X��SǻΦ��'5BTg�
�T%Ku	N�F�I&f>#,�S����-�{�5"����h�*�n��U���3m��+�%�r�AIoa*������#���ф1�z���AŘv���SvE�/<k��-�l{�'�7T%_olc�pɎe�.۷+mӹR��x�BT}�U��(�	YL��=�z����ȶE�?kl9Ϗߌ8���ɐnpxUBUB���2ȵ;�ƓvE�>�Z�ȶ=� �T%\��K��Tʴ�J�J>폪n���_2FT[�>��RE������|��\Tq+8�gVE�/���ȶ7�;���d-���Th��b��A�mC`�\Y��uYfF� 9�HY�VcR:]4��/b0���Ȕ��Ʋ�R�����IM�,�Sl+|pC�pі62�[��՗L�J�d�.tJ�1�X8?wwJ��}�;!I�D�Ԭ�x� ��>��p�<����-��e�%�,зQ�K-9_i����먢�qU�,��;2�LL��+CEj�1ۆ��J��G52�����;�F�-��}�d[��&�gY��ln�e��N������
�E�uֵlE���Q�lE����(j�����(v1��ÒڡՒ-��=�FY"��y;�v"؏zc_\��"�߽a7d-N��y�|�g9�k�9$n�Z�����E���OC,�l=�֤n�[�2*�J�߹����"�c�d-r��������C,E����s���2�&��]-��$�ڮ����݈�#�ǖC,E���_���"�Z}�)9�Uld*��v�ha3��j;�ˉyz�&MTy���LK,4���i��NL8�qk݉�c��xw3x�R�Ŝ]�kp����mO:��pu�m&����o�}a�$[!~�<n#,ϼ�<�jɅqPg8J�`b����oaO�L���s�M�b/ݳ�䌲��?Xn���מoM���'9��f��rd�Gg���y��䅱��Ͻ`݈�"�q����~�k<��G]Z�K�ג:��_~�>Y������lE���E��߳��؋R������&��i�͹��Ȍ����>�ݒ������5u#2kdƮ�GQ���R�8V��EUP��\@݈�#������^>�Z���3w�W��'SDIK���<��[|�jH�!j7�<�ݒ-���k��d�a�޵vB���,d�*�� ��L����"�k��-U�Z�j7�tx�sT�z�s�Sv"؏�;�!�fA�]��3=mê��ɜ��qYb>����d-�ߞ�#v"؋���!��>���\�ҙ"-�HV�⪀oi-$��/߹v�[����8y{�u�����O����hi?�]�\Y��,�Z�m��}�is�;m%��-#�i/����.�㙡�2ݸ������m.�tV�^ޒ�Kx�VsO�K9$F,��IoG��#^��m���D�l�mb?~B]�h̲7�oKۤ���;�:4HPS�E�j�%�X�ٵ�9U�N��;���lh[����|N�~����rp������D${����l^�oş�h��A��j+�шH�g�;:~����1,���-I
�%�H[9ތ�1!}�bB\F�+�w��r`�b�8�ӱ�\wr(9c��/l�����4%�dBF��bG<|m��A�Q�5�H��6ƅ��"3�lhK���*�}��������&g���щd�ƅ��DZ�=���'ؙڕ�#-L�$n��HK:v��p�������[>wle�V]ݵ�\K�a�U��V뙹y4r�]z��K��(͈V2����L�XÝ��',{:ak��*xBy90幆�Q��`���)�c&�3�e�%b! �z�F/�/�:6�g8�p��_����^߼�_4�Lхy
�:UwW��gwI�!,�"=�lh��ln̙QS�qn\WK6�2��
?~�_Ղ��_x���6���mE�8��䏃B�^�H�~��m�!n�4oS���ɉ�8b=���J�l�ط��bB\G���9�����g9�Z�����hH�zƅ���H�۱#���'2\�.�1!n�,hOEk%Gv�֒�Rra�Kv�����>"���vWKb���y�Փ�9�Xb�52U�țV]LiB���Ev�a���4�X#;J�z�X9���lͅ��f�������A���.Ӵ��na		|��H���"���ʪBG�!�4f��B���ʍ�jؑ���U@K���!n�4%�2UR�m=}�3���r�È[��[��*��	b61#_6ȫ�.���.�C.�NU$��>�*���b�=�{Z����bޝ;w��p�o2H�K|ȅ'�~!e�S]RƽiM����*����B�et�$/|l�#�}�;eٗ�,�%1�R(9lV��S����}�"�Fvؑ�j�,HZ��Ź̓o��3�Ü�M���*ĉc��KWﳍ����5V����G�>����2Hd&ZH�$-��XЖu�
�&~~�!-G�����ppUv�Ö�$ ڪ~��ď�;cB[��-
�UUL�=,h�_�/E�v�rL�$o߮ą��Z��+$v60���V��<�$����~���$/��hK?2!a���A�g	�K1r�!I�pJ�̯1d��#����߉�bB�뒵T9���G��^v�e�f+1	�祟�_�T�����!~���`1}��n��#��f^�ӎU���U�3�6�d+���D���n�p��H�~�;,yxGk-cP��6Ƅ�ð�$-��ƅE-��
���yn�M��	���Б�T~�8L�n\QH5.+��݊�Z�;%��������"?>~�#?{?Lx�Ɨ�q������t���bG�MV$.��bFzm�	{��з�o��Y×���|gB[�J)	g.ą����$-�{c���mv&v�dh�1d5�l�K����H���bB��D,Թ�F���NbE��>�-w�]�[�x�Z�<��e`̕���-r�-���-���մ�.M8�B%�|��CM&��v4�%�ق�伃,��Yeڳ�6�F�:9�K����"�rkd�%h��2�R�؍��gX�hBت��c0L��%ز4�1		l�k���)�`P3�۱#O��ݙ3�dBB�G�4/a�.)NK�I�V��Vɦ���gww�'�>z����F��.s��P����Х˴]�"2�)�w�N	_Q��ϬhK��P=�±#z�S��f7�,H��v*�?�E �ϼ]Z?>���	b?J��P����������.:̷�		~G���#��b�>"!#=6ƎW�vS�%�����QG�3O±!/y�	��ĄUT_�tʴ-:.��r쓆rŎp������Wt���[<��FD�Q �l���	W��W򪢿~���;����|?�9���Wfg������*lBB<J>t��1�𫘆�R|N�c�"��1J�iR��n�;tW�ي;�j���6�.R��\v�٤��-**t�s]%��津�Y�u��ۿ=^�	�t�a�W�E��ڬǖ[U<�y1�Y�(�����<�¢ʖ*��u�.;*��%��]��u���;*�&�C�;���/p�M����@J��Xb�/
"Q�u��'��B�L�ޒ�������y�{׼wX]�Rő�u��KVۑ�]�"�ep���KXbv{���\��nQU�y�cK,�&؍��%m�[��[QL����<k�QU�����:
�E@-PYjm���5�i-�dc+��1��!u�%KAIz������wj=�ε)��:\�,�L�`Zml�3v�ԭJRH롮Q�����F�Ɉ���6��ř͒T�]RgSH�t��B,���0��u1LCG�4P�-f�[{4�؅�]t��!_���,�ۉ5f�ms�dۯv۴��ɛ�B��h�Z�eeҐV7���cM�Zm����Sԓ�	��*�O*t�ry��A�vN�?��đ|�u~��Z�V$3.�͗,�۰�M)4%�4	[̡�LB]er�(ݭ��	�<�'����jH���N%.����Ow��������}lH��< 
�!-Gъ�m=}�2��YÈ[�.�(BGς�	b61#y�bU�z�㈵�˲ِH^��ƅ��"T#=6Ƅ���l_M&�8Gw.1pHE�"!#��ؐ��V��P��~�����-�K2��K�#�]�	���6��4e9��:�9{�ʯ���-	�lh_�r1s��߬i�=gL�M֑�2��z�5�ޅ�%m�#�Cō_ȈH��cG)s�Jc�Y���x��~5��5#D��S#Ǣ�R+M��m�WL�q��������u��a:��N��ju�n֢r�g-��v��+a�u�ֶ7p���C�r~ďV�_��]�_m�]{і !p�_��Ƀuyi����3��UB�J�bG�,h��Իk%�p�t�B
�sf�о���Б���?�H��1p��%�'%�\��!~�e�"A�ޒ9V�hn
F�0��YRB��~���۱#�B�u�dʉ�qɮǴ�V�z� y�x�BF���ƅ��"/���TPĪP 
UJ��$/��.�����VG�r듦��ou�5�%
BȊ+K^羲!~�2А������~��]��!#�mؐ��Wm�RePT��?Qthͫl	6[BU�FɴleL�&Ҩ�^���F��������R���R�_#��J�F�����g��=9��έ�|��ŕ�tR�EQP������?\YSwO)���~�B��Ŀ8�H!��섄"R�K,��ܢ�* �������!a��-{��|ǂrt�I�[����]�=�~�H����a��������ď�c�P�J���L�$k�� U\uӷ�$-�T��5.|h����1��QhH�a���P��ף3��#����,�X�F��R��g��cB^�"5�����)���]���aŎ��)��i��EV/]%�)�iq�m��8�U���8'Cu�DaO��^l��Q�TL&)ئ���,�Ҷ6
��ũ.]�4A�Yd���TUW�T?��|�M{��a˾E8$/ޕ��Em��M�����L�M&�j�E��,g
���KO���$o�t��~_)��l�m_�G;�e�	�eX���݉��$k7�
,HK�dB��ir'Fs������TA!}��bBߥD$o6�TR9^�n	9�r���	�x��u�c/�v$,=V����\�'�w3�8�QK�Ȅ���ȅ�_V�UR�6X��}���<�y-��g�=Yl�>��ӑ�3:J-�u��!����:�G~�K�lb�[O_x<XPQ�;�ĥVHk��J�iY1�m&8��:\�ˣ���M�<F+cI��MpJV]�^4!��d�4�!�1eX��*��!#�w�Ȅ���T!#�ydU��w2J��˲��,U@_}*!#��ؐ�eD-Ϗ�^���<9�aj�$%��ď��ؿUU"�)�J�H�~�dF��r��e�1<�b(*���v$.��1!{�4"���l���>���\���eD$j�(��+��fv�u��1��O��>N		|��$nM����紦I�"ÌF$O:ww����t��H����${yeP�ζ1Y�n��Ƀu�m����P���G�e�j����׿t�o�I ������.Љp�u�H���ƅϥDz��U ����Ȅ����ߠ䳄pŊs�B�_��?�h^�Q
�
G��#��֮�/%+��${zYbB��xlGe�;lE-���LY����(+�#щ��4-�Qy���{O����$t]I�,n�!/#c;�]�ζU�{cG=�b}�f]�S+�ힳ�U@B���/zTBF���Ą�#�b���)w��^)k����TBF3�O��
%QC��%�lbFo.Čߍ��<��8b�U��h^쨄��>��~�*!o>�G� �;s8pHKu���0xkt�6���MJ��NͲ2�.8`Us����H׿ďkći�F�Y��12�*�*����W�oną��"�{cB�ʈY��ƍ�ÄɒN`��ek�I$I�^��m�[��5V�s_��*��ŧ��7fc�v�V�����Ą���5��"��!fqmM|9,kK9B�
=��3�݉]l�{0b�2�ke�Y{�F��?1	`
�볃e5Ř��%�wP\4�6���;0O�׮��9h�Ҙi(���wm�N-Y���������d��1c�l��E���]����CN�R�8��Tv�����e�$s��t�/2Ae�BG?O��1���)R�J�܄��]5JZ�����$/��X�����3�I��89�s�DpV��6�IwYUT,E��^z����lh^�R�����H�{�$�;��+bF�K,��
�Ľ�D$g��ƅ������QE1~:/��vN���(g���/���ȈH^�{cG��aڸf<2e�B���{}v$.:�bF�,HAT�Y��i���xg�_!z��}J�M�1�M��I�)�\�}���
/��`��b=���˽s\�G��%Xx�-S�\�q�G49jjU�&:����Yf��
�Ɗ)<��[�u�ۢ3)�tkH�2�HD!��cX�K	��fm�b0�\�]�-{L�䓨��BB���4.rTBG��!y�"����d�r��ծ	j6~��EUA#��ؐ���BB��%���F��r��e�7���zm��J�H^��bB�ʈ\�s�_	��.��T�Q���y�U�W����#~���>�ϯ�)2��ǈHZ�idB���P�.f��RbiM�͈�����u	����*!pཧxreg9wu[
ވ�G1��w$8��'���H[�TBG�O�h_��D$n�=�omd�%.Lk�����>��FB�IL0�5���bE�J���cQd4]H]�.I�,jI<H�R~���{�wUj�x�!.���������i��rY�N;8��b����ωb���?��Q	�}cG��GwY\�f!QE�Rt����^�H�߮ď������:��<�p�Ws�0�%�����Db䋖o�l��8�03�w~pQ_�U]���ʈH_��K9����2�y��O%,õb��5���ʏl���D$n�AbB�[��j���$�"���!y�� !!b�ő	{Y�~�cFoƻK$��e�ۤ�!geDFўB�$����E��A9yy~��V�������:WEd�c����w{&�^��]��xK�7 ����\���L�����ۍ0��LFk���,T�,)KZɓ2�9klfͬ�sR�"jK5Ƶ%�q��T��.rw�g�󾟚��g!���L�FUI��i�����!�b�bM4#�-mr���3��A3��:ma�V���fs��`.�3���9�Z�9��3��fs��볜�m�&]9�v���j]J�k�r�j�v�e��mV�m����74��iY�C	(m��`kbۘrj�tf�`�`���p,�͢f���6�@
 �+�]!�55�k3�5�.�5�V�55�
��א���[��7���)����ft0Bvsi0�b��n a1I3#�:Ŵ�mra �K��Ru&1�P�F�*�����z�B1�v���]�4����v�d�,c��dT�%K4c,h��SK
$d�E���1��j8�!
���I`�����t�jkV�n�t�fq�E�a�C]��iX�-P��K�Bd6�4��9̀v�x�@�/B7��!#=y�a�2� m4���l�����e!��۬2���q7bK�	��0�L	JS	�h�F1������Ć�z����Uih�]R&ɉ��$GO�k{e^�{�]��xp��3�g1�fph�*����F$w�]�J�TUR��,��c�gj�,J�|�aO_l(�ߧ�}ii�L�
*RL�lV�ܗ���|E^z%�	n�!^��6�9ɂ>c��Q��K��UU��8b��ď��V$/:�� ] A#���8��z���M*�E����E����l(���UR��j��,��K�8b�dBE��]lbF�5X��|���Y� ��x� #�cB��Q	�zut�x�ʆ\��D��˦\�t��
s��XC�B����nn%�p���.Ү��M�6���Y�u#!8v�r�7
gK�l3L���M!��)�i5Ys�)���.3E^5�����	q�QX�mYpDf�TPʣ�Dv1fu���g
��סG����o��+��$u0K�b�J��\�˅�E��|$%�2!#�9cF����u�H9p�;2l]�ø��l)��8Q�;݂��lh^�QO���ڗd��+y�Ç���
bE��!{eD$/oIbG��aڸe��	���l�������MV$-u��8�z��'8'e���TBB�w�Ȅ���UUH�mؕ{O�U̙��tb�IbB�a�=SJ�Ia��5#��,��C�u�BG{;cB�^�G>�L��E�r@�zǻh�K�f���k��1nd�)�j�-����q�%R�&�=h�v�,ۗ����b
K433Y�^���}��i_4~�?���s����?/�ؐ���bG�?˳.щ�9������T^쨄���K����� ��.�����Lǒs����ī�C�n~�k����M��1����n������������w���y?=����%��o�B�Ny��wd��`QU��W�v�5_�{�����a5�I�Ĺ#�5����ҽ�%Pg�g����×�f�����&�T��b�R�j�9���Z��:@�v���=�B�(�������NV7y2a�����\��߿C�ܟ_꼲LwoY�UL�~fy���_��|����b˼�d���_�����Њ��Rn�ȭ�����&Xݫ9T�~���?s�7��)��BK�.Ɲ��1�+������Yò��(�<�_7�N,��r&WMz�����^�`W�����.1�x��o�C��%-��[�����]dq�ǅ�����p�ү��sE�ƍ��W����I��>D&� k,�r�".9pJ�C
?��=��?~�柎�ݙ�[-�G1�Ha.�D5#�+u��a~{�t	�zpѯ��d�w.a.���3����<��@�HE � �}�~/&fBe����Ҿ�ҿ~}��s<ޝ���D^+�AHER �R߿J��ʿߠꪟ�b���!%�1R�hl�U]M���������-�0��`�u�F�Ԏd�,��áX˸�[�q�I%XB2v�9LmIؙ��u����vD���-�ZWu,D,C��_�ρ�}�4�;�~��~��e�-��Q(v%�6�2]��u�	ҪжI?~�Oz�V��?�ZR�1�^d�]�YK����>������¨?�����o>��e�L̏�ߙϻpf���G�@s���mA�c��ߥw����n}�?d�)�B'���/�������/���O�Ԃ���ƫ��m�ְv��m�h���L��R˒j�y:|������}g=�U˳.���Uv� ��J�Va�u�n��+`�Xtطmۂt��#e8�Gh��̚SdKfsXV���x�iA�S�[,j^nʾ�+����۠��x��u$����	�߯}��}��\7崞K�q�V������[���5�w,�wv����b�����PUp����?I���e'�u�B�2�l����v&!�0��k�-�O�>���|�y��3��t�����\�4�u�����+weY��^�_k�ަ5w9����q����'	TYQ!a�G��l�!\��?�|�Y��#u-Ĵ�#�l/���UJ�߽+����y�A>ز�f(�����{<�U{����Gnd�v��=݃j4�Z��d�(AK�Q9D�M�h!���ߡ{��{�n�3�o��jĢ�0�&&WO=E�a�W��{�}�p����r����_Q�l7_Dsw��W��O,���d�J�������9�|h�Ri:�}~Є��/}��}��C�BX	�N�{��^>��<r��Yd�we�K��`}݅�{�ѭ]�,�yr$��iEM��|.=~�������.�Wc���Ih�F%ϼ}ϡ��*��W3���lrb�L�wet��/��aa��`Ә��?U ��������k��Ufb��c$Vۙ5��B�A�U��6��D�c�Fk�Z/Q{i��Y4��ܢS!)��i6MʁJ�oKE%�KvSB�Y�)(bf�2B�Ő�Ϩ�EQ���;]��c���
�݇�4ǒ����ҷjX�1X���ӱ'c8Tw��w�p_���П8�['��bjCu����\��>߷�sB�����;�F}���50���*������?~���o���e�a�{]^rUQ����+{�ϣ�~�!fE,�����s�{�*�u�Fg=�٘X��ר�*���M5H�m]Z�c,��r]]�w����7�9�O�v�Y̎g�i,�D�d����p�d�םm9SRp�j�J]	���К��-��	����4 qȟ&���ssk��l�쉌cq�"<�۝e�IU�]�AUn����[ΫU�Vݻ+j�vp�D�U��Ť��̈�[s���&GSgj��!�bn��U�0教�C0�m5`ɒ�Q���a.B۠�NҚ�WA��Cp��L`�b�M�"c	���ґ�&�L�B�D����f�]jQ�+c���`J��$)a�Bm�B�i`�q���:J�A����%I�zL��֬(���Z1�%Lݘ7NE��h�1�3aƶ��,P�;X�5��0��c��8�pw��T�{I�zU�L�ւ�`���A�ۖ�q�*������vC�C-ڗ�9��Y	f�)����jv1/k!�a�jJR���	$�ػ%I$�}����n�C��ea�4M�wa��Uý���n�K�����]��𼯍�\����`��^���j��a����u�v�?�X~�9�gI��!xn���7F՗��F�c�VX��n�;�|s��r[מ����;w�W9Hew=��ˎ����x'����}�.߇ߊ�4�KI�ϼ}�5,XT�B���%0�I̎%����8�-Ѥ`�Z�5���nUʭ̍�\75��Mcm������>�w��oY{͐O�,��df[��{����߶J}W�;2��c�U�f�9�pŕ.ɇ����Whf��R��t�\6�g�N.u��a�}����21C	�hj�R�� �I�����W���Fn���2��])���g�G���_�f��h�|~!x����l,]��p��zs&gB���-UIӪh(H� ��!��fiӶݘ�7q�������h��>���+�?C�^�����e�0�>=���ȑ-�i��N��F���J]�mٿn�>�,[���?���?�
T�N"ӵj[D���K��c8n��y�~��{�ag�zv[%�R�W���]>f�yo��y��Re��p^�]��=�ʽ�mo;؝��s0�����6ARv��|l�w$-g&�;H4(l����cZ�DcL0�9��en#�[.�m���z�nf�x\��x� �]S&��:N���\�Q%�\�ݮݱ��V��Xb����_�Iw�툙�q�[�}�D&���tp���V�Kg}�0\�oHs�G��53�<���%����*�c����ߡ��+�B�I�RG������!�E���h=�G�f��ȃ��|4s{��a���=�w%ٓ����vW�f�g<}5�Y��2�퇶�˶�72���j6��n3/z=~'3��a��/F���ҩ
��ˑ	e���H����uy��U��l�T�m�s�A�3&�:�M+�i�h��VV$<;����26���6t��v��G��C~z���4�~S��m��Å�G7���A������5n���Dxx!n��96��Xo�߆ڗnR=���ᬳ��E��s�߼���df\ɇ��}7�-��d�(��Ë�D���tξ�sayɦ����".�2ˉ]��8�b����6u�ߥj�3u�>ز˙��{},��@UC��,^Z����l���c�o	�������6����1eK�2e{�ʳ�����}���Ӯ�2$\xY���o��lj]���!�����v�n�j��,ݕ{�uG�2��a�$��A�!&\��������;+x~�g���0��y30��~�x^]F����fi��fF)�.a�v�\���f����,�ʘ���T�ղۄè�F������9���%�e�/����s��߿C�ޏ��o���$�p�c0�ޕ�^�,j�"^���ӇW�a?_��'��l,ߞ��d��k2KP��Պ��i��x{vW��*�l/�U���NT�v��^���H{~�����5v��yyq�a�}G��^߈n��lD�]��0瞣�+�V/���-���4��#QH��Ü�i�Uf�bF��o7�ع�#ʛ;6��GB�m�Jd�H"R���0ՙ���C�N��y6x�n��R]� ,6�$�Qb �6���}!������k������%=��zDf�ܷl�\�IV��-+#���oz��yi�$�C�����B.e�wվg>����*�f��7���=�����+x�8�F��pf��=���%���O��_|�/�P���<JĎ�l���o�=�����c����~�}��M���f֤�
���s-�����=�;�^ߡ�lK�wr�%\쉵e��F�F��j���fiXc�­�F7%��Ӏ�MV���Y���ܰ!D�L��3J��L̆��_��{�+w�/~��L�Z�e�F��}���f�w�s�Β5q\�L�oeuw��a~z����+wX�%s2���=��w�_h��?~+�VR>}��Ϥ1�Wm����^���j�o�\�%yoüעO�,�F��D�ubV���-�s�Q��ޒ����d����xL7���9E N��V�Hg�Vg=6�*^Xɇ��3�;���6��vڼ�6dw�o�!�?#�~��?J�ߺ��؇�jb��k��K��x��u	,�5�N�#�"��}ޝG>�6�㢁ucbVH�hI�;��˼�wa����,�V���������|C5�=��s�oz�rY0�a��3Jy��ÖI;Xc3�L����j;ތҵ�M��+L!�"��Q)�U>vCT��0�e$��%s���p�X��3m�2oM椚�E�u����f��k-Ӄ����N!d,�����YZےE�R�7�NBĶ-Ĳ,�Ib����@��8|�d���"Z�U�0�)Iմ��uO '���5��1��{k��-��g9�s��se�3Fi�bp��&Qbۭ��i$r���� �1�S9�s�!�J�s��jgm3��A6���:9�s��s��D��g:��k���mw`�vɓ��1�0���5�	�kv�	t��kiW@����@�(:���h�D�!�SR6��f����8@1�1e�vf�����8�
�
����;�(��6��^���bG��b͛&q	�R��B�s�$�fr��ئ1I����7Y�p�L5Ģa]M�$؂b��A��Θl�d�!IH4�� ����s�iu1�B;m+c�n�[u��@�<�Rk�����]$��a(
�S]5(��)m,�NK\�U
+�dBv��ͫYKl)0��UXgF�%(���q-����nŶab�f�L�4�z�J]��dE�l���8��L.��e�^��	P�`�B]�0�$fu�1��e�+�t�K�����`�)��!��c�O~��>O���t�����(�"��xb�W�����?/����=y&V8)�a��Q|�=���=�ӷl�ɑ����z3�|R<����ٖ�,�������_���ܩ�D��E�X˱��]��a�tuߎ��������j��.������~F��5�?ؒ��툙�q����������l/5�"�4�^V�a��[���|��� B�ۦդ�YK��d�m�Fa�Y1�9�I��T�6�`�j0�� �r��У)onįVҲ���)�IfJ;�fT�Vr��bL8�֒2m.�0��*����j����yv�.<��tu�}��Rm�f:�륔���8w�3Q��9���rLx7s&[v���"BZ,RB������[͆����S�ّ�̃��=G;�<���=���=�G���#�_���c����G�=8s�i4k��f�z��!�z���L>ؗrEw�v��x�~�*�^7����l�ŝu��v�Hh��|���������d�|V�"�ªh9B������]4�]d�]�k٫HBh�)(XK�R[R��&��6��At��Ш^�V�!?'wI<`��,Cb����p�ӻ�_s������~��>���㷗2��o�]�į|l/�W8i�iY�"y.�k�gxCw���A��>�� H^$�|>��c�7��~�g���œ�c0瞢5<&�q�a^K��2�-�e4{���Y���6�A���v!;fK���5.5v�a��sqߏ�QE����>����;������$�E
��Ab��s_�~���ߺ�Y.d2̎+���}��o6y����cp�!�Z��g}���J�}�WI��J�w30��	�\Ie�6�M2%H�ۺcPe��]�d3N���n��s����fGi� w��v8ˑ�p�^<�G9����U#7�9�����]��%��?~�U��=�����n�ɕ�)L����f}�� ��3Q�����ۻ��l���l�q�F�H_�����*bwr;����{�y�R���mΚ\6Ͷ1��A��~���Gߛ���� tw8A�q�[%��N_"7���;*���k蹢[�;b&fa�#Þ�\��\7e{�3[�.�1�����a�_ʽ��ϼ_��$��C|G���|<cA�h�~����<�ϓ�=�{n��)s%��.6V(���Rәm�j6"�X�[&�����*�)�F�A7iL�a.�RKؖ�M�2�2:B7s.��Yi����mf�:�K��UT�����c��̼]�����O�=Oa5�&�n�SM��Y��$��>�|ϳ���Q��Jv[2^<k.?��J��E�8�gk���eo�����~���������ڹ���+>Q�6\�0�洊Իv|y�s��EP/��F~��~�w$j�J���!y�^�J��՞��dX���yb/]�y݌U��V&xpKwe/3D��0�����`����9�oE��W�t&"�=�,C�!�Nb�	ʑ9��QԒ�m��e�s�$E�̱r�:�mh���Q%�hni4�J8X��%��QX�L0HHk2��֑�E�]о�}�����ސ�l37�-+2dO%�џxD;G��^�E����f�����_��l7_Ds=�}�<�e�1�������=�[��#����d]��]�ot�t��x�)����h֌�C��4��F4+�y}���bu�֬�\I�
�u$��n�w�a~�^ߡ���,�3,vdv���G��N�J϶��W��c��"fZ�g�z����}o�Æ{S�v�乖{}+���}��<j�-;2:R�tg�}	����R���Hrֶ�)��t�}E�a���9�8�`�WL�XU���g�~~�����s�%�}�~X�{Q~�ɽ��ϼ/��@����3-�}���}�=�1�8Kes��r'+�A*�@������/v���T�����Mz���=���l=_}�����2y��߰�N%����l;��5���Tv2�ߵ�!��*��-��V<�B�\J�Y6˲\V�3n���J���6�7�]�f/n��QH���o������˽Y�h�"�a����z�ߡ�ot�E�fc"����ë�37`���px�1"䅢䍈�U�
.Y��s+S�n��j,a�[����d4�m�Y��aLJ�K�LMt$�K]��/]Zq�6N�e�J1�&d��I��ћ)4��RgǞ���ҝ�̙1̆���Z�"ѶЪ��<s(X;�w��߇q�������`��1ܵ1SwR:EحY����WO���6_k����r�������U�a�lK��f��>#y��{a�s�dX���yV^^�g�J��Q��pK��7nL������o���h$�=k��k7Kh��r"ܐ���;��/�U��M۷9��^��E\]dc#im��ͱ+*�Z�Ŋ�n"�mƐz]�%vUe�iR\][:ɅY,�����K�I����U��R��Ϟ'�E�F�i9�m!��96��0��TTX�T���-G8ƤO������Eꏗ6'$��oQ�E;���$G�~}߫� -
�[s,��c!�,�b6��v�mT(�� V���V�I�,U�m�\�Q#uMJ��hb��֘�"�Aѡƭ�t�c��b��f�\[�!�4��MC%������0��v��FF��5�ҔћV�&���(��$I�h$�B3�Jn�M-y)��(��1H.n�H�ka]p�biX2�H��`�a���.�'6�CA�e
��Sd�m6ƕ�`�,�ԜVb2�i!��2�I��:�-�WQcD�ٱ�-�ٻ7	1�[7L�(�1L�O�]d<RyGgr����
=EUQ��k���M��vEjF�;k�[2��31)��(�Ʈ�I�R�i���0��C��̔�J}��xx�y,f�4s6SY��ޏ/|�{����h]�G�%�"f�H_�${�݇��3�(�,y0���9�+������B��ѓ�ú�(;��A��~�G{a���l�wN�Y=��KV�v�#�B�1�nP�X�.��7���������%�3�3�lk�.ZE�!(��"-[��.u���Qu�C7��%�&c��,����)�U2���d'�4��t��y���.�RN�eovV/���.k�7Q�Zvb�R�+��+��{a���Y��Ͽ~sГ3�K���=��2�N��2��ա	]�!v;�������^_������y���"J�Nl�]2e�$/��=���_������X|��=�霁�{a��}5˩�]�k>�����UY@Wߙ{������e�$ǏQUE-�����������V�#k�Տ2����	���5�ЋpW.���2"U��X�wݮ��3ߓ�>}�{�:M�CbY�K��_��D�?��A��ޓ�%��Va��?UP#�;��#�?C�����<�wP���6ϡ��(7�5|/˙��C}�̙�0�J��7zJg˩��oM�`�i��(F�nn�`mƤ*c?�m�M]���������e;c��+-���4]�֩f4.�e1	Dz�I�$�X���zYmfK�i�i��ԩ������w2B����)e�nf,?w�?���_�E�?�3�ԉ6�	H3^痿��a��\�i�)d�#Pn�ʲ�A\��.�Q�~!��W�9�J��p�`o�������ޏ���ȱYi2�=��Ͼ�����pK��6�,˧Vsv���f�ˆ��z'N��o$���Fm�7�.;�j��D��Ƈ8��ߓ��矣���o>��f</0Rb�b�%ږ�[��e�YqѤ+6��82�e�jSy���7f��e-]`�p�Tv�j$'wpwÃ���M&եcH�;�dr_oH}�ʽ�n��{iE�cɄW3k�w����+�6~�����A��8�L.����˂���=�C1st̗W"�E��H��^�G����N�e�˼��u��`ar[e����؅�.`�W15������ߡ��^��n�ɘఏ.�ld���I=��y�n������D�Լ�s�o|�\NH���jd̕1#�	�2�8��Z�Y��p�:0�Xd����':t�Mk%rA�5)JU0�Mj%�8sn1�j&d�iF�2�6\&���%UG!V�+�
�:����QU�{IY��_�����.�Vb�R�/Q�t�������߇���d�����9��{�+���=�y2��w���=F�HY�"R��Br�11�"�������V���!<���� ˘v�HJ�BŴ\.���F�l3�Ws�]Lyy��W�I_p�/�Q��g��\h��2f�����Nw�\�&�-ETR�8�դ�5-8�]�u޾��3W5#��Տ2��⪎��u߻+W���y���*���a��ub�R�3I�1I��f��=~>��p�����~}y���K�`�L��-2J�v��Yxo�5p�3v~*���~����{Z��(HY�?N����sCW��~��e�2�w�����!�3Q���M�R˴���}���ў᰺���❦�BYA�RS0��M�mֽ.مr$�Ur�s��U��Z�R�Q�aؘVVX]�eR�4�X�Q�`���đ!H��;�����j^p�1��ª�0^�W՜>�C�p��xyx�[,����ak+i	e6�Y(c��;��/vg����̻�R:D��]�"��1�!�}+ٲ�����,WV2�9�Ͼ��ƺ��9���<Y�N���9�:���텞��fg�!,8�O��'�߷�h������Z�̭�!�^ґ�-Z?�����,��t�h�{��>���#��ޥ�3x���L:�`M�F��L��������#���)Ry4�gT�+��q�SG�����a�b��e/-uW��]Ĉ��8w����ej�ў�繬���$���_u�����.n����Y�߇���Hf�G�a{�]�,��2��g�l/����y|k/~�Z���b�L�O�Ͽ�W�!��d$"9G � ��Ee��z}��V�Hf�tJ���BM�ê��k�����x��᰿l3w�]���1�3/�Sy�l����q�ŵ,˅VPQ�ジC����Ù�8�`�Jf�^�!ο���^[��8�U��WI�
~�˞��>��!���}q,^D������_��ȭݫiۊ��jB1�
���.~��*�|C5�\7����O�q���8N[�Mݒ�%���߉X}�^����3�oTh��3�y��_{+����� ?�#�{�c̼�hXw������W_	���� ;AepX�"͓i����Xp�s
��Rw'T�u:�1��[�Y){.a�}�Ц3���!��=t����&���W+����:��G8�UY����,NսI؇��`���\�fs��i$�N�)JC�.)L&!��6ҹ�s�v��v��\�Ύ�-��]��39���g8\g9ְK���JWZ�	��Zo���;Ͷs��v s��l�Vf慷\�̳I$aDf�l�Y��t쬂����Af��4�E�n�3q-���kLb��(�nmI����Ę6&ĥ�w-bͶi�9f�h��а�e�Yk�;V�%�K���T-
y/����ѥ��W��2�aL�3	sU�i�$ё0�G`�İ�s��f�F�
b	�0R�V�0���^B]FR�LNK����f�D�0�60ۜ�]Cg5�{��WIi�Cf��-�l���a���!Ha��,��)Cv�]����kek` �F�R1Epf��,�Jö�ŀ1�%Yr=���I�%3J�]����R�d6�Jޙ�Jl[i���^�$���1pJˍ4*� �F0ݷX�؍Ve�Uf�������qHR1��Q1H@��{y(�ʇR��ة��;����Q�z��JʨT# tF��%Yq>���r�P�wa���Vn���9[�>���K%Yxo�5p�	<���-�N�D�Ȇ�%��n�9��{6���>y�|R���KN�g�`B�'����A��/�|�}��|3&��Kq!~��N�P���c�����f�u{IH;��o�Wl/�U�p��x�2e����w����F[r1�!17ƜQ˲F�Z�����e�˦��ukq�e�5J�0�:Zu���1!��Vm���u�
X.��m׉,!�SqcЛ\F	�c�};����W�1�vay���텊�v[��:Β�%���>����|�k���|l���*)�]�ƕK�wc��ue��=G�}+~���f{{��	r�ewvT��<������y��C�+x�պ:��п=G��߾��f<1�Lŕ�v��݇�f�sv�N2<v����^��nȪH�n�NR�d�h�$�]�>�t����i�͖��|샓��H�0��W����܆e����WiACB"��[-�=b:�Ͳ���N�s
�)�Ԅ�l�Q<��|��7矊E��	��:����_:��k�g7L�ur&dx{����3vV{a{���9�ff"�0����=����fo7��]<��l�f��9�������x��Ѩ��o+�l=�o<�7C�!.�"BSLl�[�{�Ý����Z���0P��+LHa-�F2;�yx�Y�����EU7���o��=f7s�7��t�+Ii�F#6!�:� -{үy�����s����[N��0�_�f}+~?J���]�<����UQT�o�{�F������}�����̓0իDz�-�v�W�ܕ ��ĒEڸ���;�%{{߷�6Yyly����v;��݅�-aW~f�Uf�?����S̙yq����UU3��?/��8o��[ߛ�Sʝ��eo�Һq��PU~�!�������ٓ3��/�Uo��W~=��z������O��5v�e�f���,��d�J��e���`�����ߝ��z�=�	>���Gs-�i�";%8KE�KXy{Y�~��=_�o�����	��%���� �_DoOпߡu��T��L��稳�C��f����Ԏ��8Yy���a�?���*�T*�!8��8@��l���-v�����-Z���X�+��	�fǷ���m06��#`P�i:jC�S��Ch�G\Mm�,�Qі����Ga&uXLY��81K��qˤA�QE`��b�p��ˋ���~{��ѐ؀�lL*�jĔcE�[�������_Qg�Ͼ��'9��̶��"�n�����>���<�a�}�8�f,J�Y�z*��a{����3�tX�Xe������}��n�3W9�Q��o�0��=��?B����~� �<���\g��IJoq���fhSBj�1b�.���C>5�w�{���3%�(�!J�uԮj��q��׵-`��(s�j��V�e���Z	��.� �Fm �ִJ|�;�
,�h�s��Yk��O3Qޝ�5�3���}�K���3]=���W���k՛ϵ�K`�6P������\����G��{�����������*�݇7�k�fK�̙]?O��~�U|�D�VHi��h�ƈ�.FY��t��}����)�f�"��#�n�]��P�M��#=����7����ߢ�y��t����Ӱ*�ª��g{%Y�Qf��_>�N(��y[핇_��K~?C��Ͽ
L��&a���8w��z�oa~��(�/q���R���W��]3Lh�GWN%q$�f�|���Xy��k��<�M�$����nҤW��i���ӟ�!�gMgƳ��{S��7�a&�J��ʳ�/��w�c�Ħ"�����w�Ɍ�-���-h5��W�EZ��~�s���qݼ���7ax��oa� [��3���E�x�᫿�����(cqƝݐc�P�����3�����w��}��8%vB;q��mƥ��	�W=����Gl/^��ߍN��2�̭��a��g��p��D;�[O�Y�����QK7�7�<,῎�n���??�ϻ����~�J�؋d�dV��ɝ3^�`ʪ���1�b��ÃXCM2A�A�V�ܺ��et �!�5њei!\U H�ٷdz�	�d��˒7]�J�%�g%dػ����e�B�ڮ�C;�z'rb�YN����"�V�#���j�M��開�.�ώ쯳�9텟����Rc��1�<�\b(h.�eŇ��#㝅����9����b��L�gl1}�=������G�c�3�ef}k:#l9�l���ڑ�{vWW�̳��UU���9�{�ǖ[��o;�=�����lXvFkס��]F��,��ӿ}+sa{��$Ǿ9���4ύ�k"ծY�����q�1�I4��,bΒn�Lli�'+�))P�PU����nƷ�VJ�:U����u��'Ruj�y��۵ww��*tCՑ�w/#�
���׋3KV��m�No��G�WА#Č��'R&��*��oS��.p�i珗����Q���xxU��̥ʎR�@�R�g��5����F�*��1�cY��CmX�P���0���v
�P�Z�+eV�[v��j�HZAmUm[�.9���MD���a�4�V9��ڔl�F#f5׳�{⵩Һ�]l�l�c���������u#L)	6l�ٓql�DD,�gHt���o�|��ѻv�6���Q�Mp�M
�F��C2���R�=�HF�'3v� �i��$k�t�f��Iv�%��`f�	���gH�hHQƒ�f,G<�WK��I���E앛i��mU��Un'�Hj$����]j��R�x�]�V��'��=��*#8�V�5�EXJv�Q"�3f�`�Ii�Fe4�bD���,%��:[��;�߂����kK��u�Ywup��������W��ej����}�BX�������>�V�[�ߵ�j�R��/0߶�pG�l/���b�f[%�Z�k9������^ymI�f�E����4X�P#����Y�������B�����s�ߏҹ�ض��>q��X�u��۶c���}+9��_�a��i��I�p�+����_���{g����Zv\x�fI����>�~�����$;/"�c3|l;ϥ{����˚���=O/-߉��翳�c,��ă���4��*iB�^�z_�o����v��y�i�3v�Yq/��N�xL�^�B���5bK�G�~b��1{enl�P�t���0���`o���?/��Ff�S,�K��1������^Xk�k�.�^K/&<7�+��+=F��/y��I�%�<��פ>��y�J�,QЙ�8@��w\;އ>9y��f�ju&I1eۧ!����Ym�yZ�k;�a�l�saÛ�Ӳf��rY�����=��kr�p��xw^�9�[񲽆�3���B9pC����8�F��,��?D�w�rM4ЖQT�T-0;:`��nv�RDҫ2���0�ٚ6c��Z¦Fb��\Cs�6�ku�!���Gt���4r[Ό���Lkyq��1�	%�IqLR𪡅{gK9��Tn̏�8{`)�w�`\�5�a��=�m�9�zgQ��7�ڴtXch�i���Dj�㱊܃���Ë�3��Xy��n�p��91�0��ϡg��l=ϵ��u̙�g�һ��?�������Yn&dx%�_�s�!��݆o5'�T��*�u�7-,qۊ4��"��!		YuvEf��G�rW�6����,x�����1[R�#�v��ɓZ8lTf���5c+ �c)ט�nfİ���MI��a�� �kl��WWIEnYq�����Q�>���PU3������zPW�����,����Ú�g�|���e�^G��6W8}��g��-�:���o7t�y��݇�
�?C��>ؿ^L�t����ҿP�g�ƢB9	^��a�W�����}�ߝ>��?B�N��M��W�wjn:�R,�q�.���;��ސ���=��i�q��y�5��QҰ�>�p��^�����	�y�٘{�ü/�B����C���3����F�7��_{5��ސ�7�C�4+���+�l?P?R�ҵ�ԩ�76WQ�1a�=��9��o啻��ɘ�&�B���դ]ڍ]Y��6W>�k�퇰z|w-̨[G�Hg;+ٲ��k����F8K���^��� 0
���U!U�0
!��[�!���P��.���g7af3����p羋T�O.c����o��
"rT��M%wc-�A�um�]�����>��3C�7�a��x���a�0"�U��{�3�����U�k����̏ٓ�<�~��\ϡ�p�{��3w�܍)u���.:��k�Y�-�n�QFbǇ�
+�Xs�!���O�K+������"Q` �Uvb�ʷ�[4���]��6�#�M�)�b%��R����A1]
KR���q�װ���6Z(�m4Ml.��1,)�YE2�,�W����ﾝ�h�X\̃gߓ�}���b;-�6��<���NHYnݝ�W�����7j8Gx���]�!�Ԋ�wNIr��῞���,��=�!~�d�dɖ�;=�è�����6���3$�H��]5���=��_��>���W���u��f��ᯞ�z�	cŔ�/0�vR��d��;`/iXq���#u����ߓ���[�!��3��W��QJX���7ιU���4k�[s��Z1$������
VҋR��%.i
]i	��a=��wpy��䎘Q�v3.}�݅��oHo�U���A٘�s.a�t�s�a�l�oпpړ���4����!�"�af��z-��.Sx&a�z����ᮽ�a~ӯ��yr# ����:xR-�G\D���彍�`}G��N/�B����8��9v�� ��]�tIwJ\8|k�o���_������I-���%P(EUS����\5���r�;O/0���J�{<�V�H{�lD��'�9,�.u��a���;�k���WE����Ԛ��a��"��+ٳj|����������.��%�-�Ll ��q�r����C8����ˆ�8���c&+%�x{�Q�;\�w�9�_k��ӻY\݅���]u
&!'U��4�.6h�>���KCm�K��Xi�ͤN;a�T�%J+Ja�h�6¢�P�I���KL�2���n-�-�Y�����٬���VJ�-ӭ#h^��!��� �#��O�E�����y9L��ɭi��O[�Y�s"�{����"w6D|�|J�klu�1ºX�K,.�..f%\*-�J�ۮ�&d�p�WVm9)����ۜXΚ�nںt��-���Յ@F���,R:��/.E_���"+��譃�=��t�����M���B�u�R�.�� 9�s�k�馚3Fh�p��&�Kn�LM$�d`�;M�nh`�vδLuq��jec6�9��(g9�s��s���ذ1���rL����:Qji�gZ̉I��;��!���3�R쵷L6��Z꘩r��Yq�T۰SS!QY����m�����V��=v0b�hlڳ�
�Q6ٲ�0Gk&��Q�ͱ�Y�-r�l��k���,�,�ѓGf�&�b�mIS���B�tdKI�	E%.�t��Q)U��Q!JR�n�͙�M\n6[*�h�C	��;K�(��J`@�%�#k6�b�-�J"$�VV3�%)�3��;`D�Q1$�-Ƅ8m+c-����arV궹l��#`
��p�M�@��ѣJ5���!a�
�Y2�U,�2W���i4�DITRS6��R�֎��,4�b��Hǃ;Uv��-�bW�)N��K�u540���-��1D�!Ham��i�4��$���O���J�D�O
Ghz�uW���S��P��������}�;ynfE������ߡÛ�Ւ,�c������F;{
�3K���b�w+�m�������,��_k#�c1��f��2��%���Ǉ￯o^�����^n�;��whʃ���}���p�{_�޶��f,xp��Y�H|�����u߳�C�yZ�}�,~~��*�R'��یo"��%�UM�v��J�cWLGQ�ΛڮD�l�˳���e+H�k�d����S�)!����b`l���Z�l���$kG�X���C%Z�L�]֕�A<�!�H~ǟ�����R�ǄW����ފ8��r�8J�vA�)".Զ��U��Y��oH_��!�?QT^,C�iK.�j��-�+���/�o��{�s�{Ln#ǆ�z�0�5o��l9㆝L˔�.��C��*��������4�W��y��z��Cx=U�6�_Fu"��\ǘ}���$��,��$���!�pe��]�8o�U|�}��9��vbπ�)�uD�nX��$�w�k4W��:m��;M�u�#��yE�K1
��38.`��Rq�d��L�6b�v;��yj菹�ǿ� f���~~�Y��xd�ߏ���Y����+3��o#ˍB{�Q}�Z�����}��Km^����n[��}���<Wy��~O��{�c����T�Jm��Vһv]�}�>���֜��'Z�L���\�$�i;f�!�rW���������s��#=O.�Y��{����>���B��ސ�}��]K"��ܖs��W�����~��,��}�x�Į�������C�~f{a�_;:�n�V,n��zA��*һc�a6º�}�O=���W��jަ�K�x;�L��-"���B�&��ޕ�v�g�{�=���nXQԷ�}��z�������јu��a��>����EUAE^�J����6���[�{�a߾���QUTa��0Ῐ��*��������߷��kil��慰����Ͻ9�=�!y�z��&+���B㊢.
]��P���}�8��a��0���ň�ŏz�>�|��s�Z�t�ݷ.�n��9+��nՙ��FD��f,=��Ͼ��z��T
�>O�%��F�2�U*[SL]��l���
(�:��v䄎HL�B�Ē�SKG�L&ٌ�2-)!6�����&��N
蛝0�M��hm�ƈ�:�^	WH�3��� Q����샐�2��g7`���,�[�m
�h��lfFo|t3�a��^.��$�%�����Ղ�Ywln���Fa�{~��l9������>~�GL������W�;//V�xn�V}�7j=����GR.��n��B����u����_��KAًo�� k�dp��r@���U�ݪ��H�P�=ӿ}+��3��7��e<WB�(ݎ�W�
;R=w\�]6��\R\�̤&d��E��1��b[�B����1�?C�ߞcԐ��H��W-"��a��9�[͇�f�qx��ys�j{�*��n��[�u�L��8����]	���P�E����ivIs%��0�U��w��~�{�Zs_P��2�2��6�-�-'n��zl���b^���Q=���7�����g��%�ɗd�2e��i܁c�V�Xyo�߻,�w����eԲ"�Res�PYU@N��#�l7�=[��;�^%wXyt�\��yo��6��w��\xb�g�(��C�vU��o�pY�[�N^]��1a�=G� �y�z�L���"��&	y,	���������[��sy��M�/2�&!%c"hE�Z�R����Vq��߈{{9��7s-������9Ӱ��[�B�7z��Yb��׾6_|�T�TP��ZSMX0�ꎵW�w�����;�.�V�,!��e^r�p_�)oO��ϿC��qH]B�~�'�$��h$�X���<7c�X������a�<4��nK2�0�&8ӹ-�bB����]�p����!��ϴ���ԳJHxX>�˷���k�s�؈�%�f[��|ϻ�V{en�B��r�yr��7�q���J-Uz�Tđ_8*)�ƍ%0��JwpJI��9�� � �ʏ2��sڛ��tU��
������޺�(�X8��9��L9Ҏ�۫NaJX��f�u����6�ۦ34-�i�̈́+�M��C]��!rLg9�jI�e#���0�e	3���A������q|}�[���t�=i�g��Mf�&ݸ�Al�h��Ӌ:�sa�4���bm�niPJ+��J"[�!ϻ+sa�g{\Ԏ�yxZ�c�~��G~�?#��7��U@�~蟄z��%�y����;��߾!��/�s�h����7�~ ޟ�=��~��x �o����y��U�0�&���y�l�m��m�@��2
A��d��<{�s��T��`U�|6Ͷ�m��lUT�8���>��9r�D�9p��ǐ���E�u]���ï�@���'MĨ�:򊋧7*��5I�RsQ_�%A��f v҉���H��BVbC0$N͙*��J)�9�Ȓ<iIUE,�R��s���t]'���|����Jyѷ���oON����7��Oy��u�_�{�?�_�����z�>������F�����������&�m��Tv;d�y׽UT��'���������O���U)��/'ץUJ�p�����o�>/��/Н�NO������/e��[���eUJzR��}��Z�irV>+뷟MF>9wO��9���"�:��t^;����c<s߯�v굳f?��*�Nﵾ�v�����iZ4%�"a�Xh�2�4�ha�4kF�f�h�h�Y2ѓXbу#��щ��U0�Z4�ѩF�(a�4&�.@�j��&M44j�C#I��єѩa�Z+FDɥX5�F�є�j��FSCUa��)����Y,2�SCRh�22�F�a�SCJ�A��2����a�Hhҥ��L5Dh`�F�-�XeQ�Șh�F�a����1SKCQ�a�42&�T45Uh�F�d`��Q���9�'!��5U��U��X12���#*��Y�#CEhbVFR0iI��45F��F2dh�ɡ�#Q`��M21�23C43RƆ43#0cRƆY�ʭTd�SC)��H�`��RQ�h�W��~�[�nKߧO����</����J����Wl��=O-�y~w����{��Bw=���_[���?/��>�eUR�>�]����ݟ�?�?�uo�|n�j���t���c+���-�/���~����}R��=����:l�o�����/G������wMO�(*}+�U)���r|y��Z��.r��z?Q���u�J�u�槯!N���lפ�7w�N޸�*q�NIת�Nn_�:���.�雚�rv�q�~���UUJq����1�:�G��TD����J������������|+�s�N��C��7ԾO��~z������+�
���
��~3�L��O������O���^��O���-��B��R��(��X��}|����/,��_��q����t�U)��Oj{��Ϛ���9�s���]�@���\w������}w�����O�b~.��]>T��O���*�S�^���}_���w\_5��u���}�9�>�^���<��]��B@S��d