BZh91AY&SYzuu|�n_�rqg����ߠ����a�� <@   ����J ѐ�  �  e� �m�{�@�@U� : � �   � `    Р ��@%A          (      �  �)嵙��FZѶ�Z�m�L��f2ͬZ���j�R� �  �|>| �=����.c��;��wbPZw:Qvr�C��gA��� 6������ݔ���є�>�{�� �zUZ@ h`4  ��� @]�΁��� �
 �w ��J�����6�٠tQ� �U�}�� ���@ 9P��@H�Z�QZ]�v�� ;d6 ���B�	p��  Y�.��(wv� l7s ΰ��@M��@ U �` ݀�@� �P��>���&�e��0 8�@��c� ֻ��4� M`��;4 WgpCA�C�{d�<��і  ����p ���v ۹�hn��H� &� )A@� �`\*v�� 6��i� ���hh�( 6u������A 
 Su���p=�,@ YlP�� �0� *��� �w 4ԃ@ԍ ͑� "DU<=Ȝ^jns�h4 B����A��g8 ���t��J t�ã�P9
RD������  ��lH:�BP� w` � t;�@�3` ��:�"                 ��?	JR��4�M������J���ɣ� �C  US���F�U"M0CɀFL#L&�~�T	*�F�L&C F�	���S�T&�UU0� F� L � &��DhMi�)�O4�ed#�yM�������0��?�O�NQ�ݩ���}�t<=�]����  w�XY�����I$ ��% ~� H \������5I  h�����_������̲�9�<~�����~��?�����>����9��_��ݯҿ4?jB�8I Y����=������I$ W�,��~�`�~*��������V�+�e�$�@ ��³���o�?����k?��� �H ۯ����I]v���1?Ŕ �����"��*�YMP�)��mFy��u-��e�P�t=��h|N�g=��n^�;����=�7q�7r�8�;���N;���|wӘ�'���}���<s�Klb҃(+*�Q�*�b�AB<5��3(�gC��M̺�{�Za�㍢ʘ!�U,r,]deYw.�eRR�IR�n��si���V&k.e�c�-�6V�v$n��=xl�j�[��S�YD;TC�Y]��!M$.�C�D�m�\C�A`������%�%����Ns���%p����wͼ½�bk��Z.`�e��e�ͽ�h7�t�a��ːl�_
%õF��wP��i��K��M�X��P�R���;ۺ�+2�e��=�eIi6�j�ɻ�]��5ૢ���іt�˻�#CKw�vgq�U�2RCI��v���Y:6���o�{k�a���|oZ�J6Ŵ���ꃦ�LHo(�U�S.�]QU�L�T�)i��P��BC�05����D���r�B�F\������Ld�}2�Dː�!�����Hr������5����̻H��흘J�*ʗ�e&���eJB�g��s��3�_��f]��\�<n��m��8N]����Al+�@Y��*�
"���Cڤ��e��cuD!׌U��t��Qj�*��XwT�FZK��㫢[;u�(A�!�SG��C��q�AY��ީbǬ���K��j�L���Cާ��']�l
��lh����l���(iF-*5(*��!T��A��#L�h��u[PFWh��mޘ&]X1��q�&����Q�b�3dDjF�W�g�����b[l�[ �������zo���5m1aM"��.���d���%�ʕV��LM S��'�[���S�"�"�O������<c���R��f�\��yNs�y͗;�>���q���gk�ږ7bmŜ��v\^�#U�|�%�����y��H����]tD�#��XԵ�C_Gs��J2�J"���_Uy�:����#�zv���q漍�VUl�k���&dn[�u;����c���vtu�>�&�����ϖ���Ǎ���υ��3��;&|	Ww:��=V�n�"����{s��ƭ��9yr�D�-�b�'������Ѯ4c��ʰ_&���t 	�  L�EU��hB�d��i�)�@��"�$&j���A9<�,&8�o�N�>����Vq9sռ�:�O��F��0剭`�z���f�-N-�v�ަ6f�}�)Y��v�c�Z���:��\������pb��\�1����6�%L���Ʃ�5׳��o��T�V��k����8�M�C�%�^NL��]K��� ��  L�d 12  LL� 5R  �̀ ��t�#�㈹_��p ��Ʋ�
6fYj�^�e��)S��GyR�`���;:�Z�h�y�%Ե�%�]u,��ϩdf�D#g��(��иPh�Fv��������>����Z���37��1+Y�U��Z��k�{ʽS��Sy=�j��Y_[7���_]}�z�1��Jg5��&&v�Kր���`�R�r�Ĥq�)uU)`)J
HJ��!8%�R�.���P$m�W,�>�D����DI�:�&e�3���z�g�<>%/s�HԱN-υ����r�5�X�G&ҧ����-����5Y���kS;s�ڻ�O�s�JR��T�75ķ�\2X�z"5���y�)�BηZ{�=���3�����YWs=J�it�Z]jF:��S{)R��2���`Ѣ
���F���T���w��1�Lvi���N�SLqщ[]���_E)�L�ӎ�%y�m<�����>�{)�7j^�t}�B�YlYl-��-�m��L
Ue*�H�)��-�W�}q�$=Υ)vy���Iu��wy�u/)�������v�tc�k<�i2�Q]v�}��Z^jX��}u-Zܤ�g�8�y�-ާ�1-S��:�%皖�pR\y�<�'�k�[�Nޱ���u=޸Ʃ���&�<�ľ�bu��%�<�]j��S��Ƽ�ױ>[Z���8�1�̖O��rR��v�@`�y�c)9,������؛k�ǝXe[��0�QP� > -Ӱ�t����s}����Y��c6&T���M�d�3n>զ
�����d�,ً �fRJU<�w)=�gkz��1�ǲ��=�<�-}@Μ��5#v&�_�ּ�S�S�cZ��"Z����"e�<���O{�s�>�[�O�r1�8��v'��0q��3^k��J�'��R��|��>���'�w���n��O�q�^���������;X�R���]�_W���1�"I�����.�~�y�\���#�%־�8�n�ĩJΩ�D}����81���j��L���o{�r�km*�7��f(�7&^��B	�(��m�0��
�8����;���{��s-�T�މ�w�Ry�^#�y�z��������n�#2g�/�R�����{m�F��$ A����|R��JF)@�҈����G7��z�:Ru��빮8��7��e��_y���1q�J��LUk�}즫c�޼:�q�b%��۔ž�dN9�לk�=�5߭��<d�'�k�[V9ؙ�8�R4{bi���	���� 4Kϓ�8�G�9ؚq��s��by���k5��܊1b�{�2ה�R�EdN��rݼ��_��'��.&�Zǔ�T���ۑ��r����=h�;�ya؜{ݯ)�|��&U���M]qj��8���tf��ˌj6�r�R�Tf*u���QY��؟w�}�R�r&���9(�^c�䭵�ך���}���ϱA��&f��?��]I�T5vp�A�6�n|�q�w�גs����n�n6��5����'�p�T�-6���Kwm:�璧��&G/�ZU<�{�S()�ɧ\���3���|�T�N�)��<�r�QW6ǚ��ծ�iL}���"�}>�q�n�*�O�����}-J]�J\ff�[߱�8��qO����9]�T���jcUk�2IN)5�::dv��Fru.5�%ltqO����yǗl��R�(�Uܯ��-,s*�.Wgk�-������T�Lwmb��:��M����k'k�J"�6�iMku��۬Hť+�����)�Ե/��ؑol[�v�u9�q.�1�q�>)N�'�R��F����YZ�Ԕ�vy����\��R먮1���.�B���Z���rMv�iBמ�9��٧M�J^WzV�W�ʝr�޾�A�n�+(����K�v��(��$��7�I�N̅���s��͑x�dÐ�T*Af@�Qɵ��2�<ԫbz�T�Zʹ�_��/���N7��MU�*9�X���]�݉����>�NDۏ���-n��K�$s(������m�J�ž�g�Jrc�[�U�^vͩw��ֆϚ���� D��u@���zd���RnfJԦ�/�ʛ����;�#Q/��m�W�<�v1�=���+����bRԶ�z����^����R�Fg��;�.n�۔�rJA�.94�R,�gf��8�^r�J\K�N;©�j��U�uR�3q�\�)�5n�*;��s������g*3�)N�Ls�yjbR�.�O:��q�j'Z�<��X��:֣vm���[͘թ`��T�	}�zsn�UcZ�%[u��1�8d��t��31�M鈘��~ n >T�T.���j�W��+�q.�VƱK��c�q��H���J��=���uo���uV WWV-+XLM�K&$ �őɰpHૺ�)J��"@)�#�u ��,Lą	}�?G���ҶܿUW+*]b�c(%�lE���c�OyY�)ݚ��Me��J둎%��1���s�޳����tc|���������P`E��`����0�EP�0Q�94r4elW�!JE�̝�ʛl�b)y=�W`�Z&9���_J�s�u�e�~ќ�vu��w�5�F�{i�nv�,v~w���EOX�����+�:��2&�W'-�T_��Z��$�yʨ���ԙW��)���=��n��t�˘]E:�/	�Vv	��`��-Q®����5��r���]c�y�։������<�ڋ}�G�d+ q�@�L�֐�ߴ���3{�v8����U��J�\���T�y�ʚq.�ʘ��W��H��K_*��}�-��e�{�1�w8ʋ��?Lu���R�����e̼bR��SIJRvn��JR5s`��)P��JR�
�oQcz�3�b 3�cc`jJH \�ͤ�LʦB㊪���m2�$4���[�}�pu@�)r� FMըJ@K.�"D�]�`��]��-)JGn�-)JR��ե �I]�����A`$Z�d�����Kl��:�1�'ٕ����R�s�U�ͬT.[�l�.�?a;���Gڤg�NR�1S1ڞGS�UByY97�f�,b�_+�Sic�������]}iu���U�b�ܶ���X��ݮV��s]W:�����}��R�|�
��)W��ˬ'�}�>�9߶��#jdh�����1)�U�k'�6V�2������ZA��	k����w^��q&m����±�����98>t��g\�:�:)�Zǌ����w�U�'�>kQ�[֋0�7�º�eB�lEͩ7$�g�g"}������q�;Dq���u��)�\�V8�=HkX�Z���%��\J7͕V���}"�ZVw���)�3s��u�1N��˩}.��9)�7��}��3<��[��)6�\c��9{��1L�[yN�g0ְR�L�x����\���'aY/*g۾����M�g��Nl[�KZ��"�8�S�����eDD���X�ye���D*��U�a
�@YuR2�
�v�U��2���.��8��YPY�H)��!ԅ�Qi���E�%	�ْ�&���˶q���p�I|�WeKMCVZ��i,�a�Qc'Oj��i����!ƘTC�D�wTW��K�ZPP3�)�h&��W(��*+���5R�#I��i4�I,����
*���P"׬�Km�Uv�]�X��v��n�,��ܧ���n;u���U������(%OXX���uXʖ2д�̸�A��Ai�UP.ŢQUQ
�!UD+�B��UQ
�%�wP��J�4� �2R5�B��RKB��)���Y
��S.z�`��h����|�F���bag�Q�([)����X��P�(�%5mKKK�
մJ�IM]X���JeP��]�]U+)���bP��.�J�Ѕ5mX�-%]�eJ*����6���c��{x�8q��whQumJ��)�v[EP�1d����������{��?��2�~������?�����DZ�(=KG�?�H���ɩݽIզܠ�6����I�I/�	��;h�΀]��H[���5��m3�ϑ��zm#J��u&�+��=��Eҁ�S�  ��wy@ӎ�B����9��W��%���u��ˉ
�#@�T�����(T}�����O���C���2$�e����t:5$�2y@`�:�C���t:z�^�W����z�^�W����:�i�%�S$||�a����`t:�ht?Vr�C�_e�Qt��C���t:�C���t:�:pD�h�a��t:�E�I=��\�b�q�YJ��t���tJ=���Ш�1��ts��h�C��=C�ٺet1��tOP�~�`t:��tJ5�t:$� �wĺE����D�pt:K�P�~���n�LA��B��z�d6� vp��Pt?P�t'L���~�?�?��z���k��u���.���"�
���C���C���m�	�П��Dt:�ht:��t;��t;�����g�߃SR C���uL�1�C���.�C�.�n�$��d=C��]2��Q�K����K�\���C����9C�Ѯ�y*�&�*�m�)�:��֤��C���t:���xI�@�p:�C���t:��$��!7�D����t:�C���t:��0�a�fC��v��:5�d�N��C�Kd~�t�%�����Ԕ�x�޺͝#^���,�˦X(�8t���GM9�B��wH�  G���t:�C�X�ڡ����M'�8o����m�Y/*�|�����&It�w��m�ݖ��0��V�.r�#YS�����w�ӭ+*J�g2����[gᴟ��>ɚ���+^�$o>k1��Y�s{���=;BS�a�ʜ�j�x�4��q�&���niA֣-:T�����yp���Vף����g +��g{Si~�M�4Z��ϝ	��6����湱i�:�p6X����"h6�&r�mJ�
�OÐY �ظ,�@zI =m��I32�䜀�I{~� ٰ����9$��$��$�   �$� {ր     �9�  [h   I$  ����z       ��ٰ  ;��fg�,��$�H$�nI�Y�r�9�8s��I$��I��Iu$�Y$��Id���C�{����m��$����� ��� ;$�I ,�@Y����d��$���n�hp��4�`4�\��e��HI$�H$�-��ޞ��I -�{ނI$�H$�m��BKm�����hpK�nfv�6_�� I$��Id��{$��o9�P  $�$�w��Phf�hp�u$��@6��[d��$�H$��rI���'�����{md�      ��32�  ��      �Z   {ޛ�      9�     �  �@        $���        ��@�$ �Z���Km�H$�Im�����f�6l� � | �@6  p�m�`����]or�9�$;t��4�g�*��{��f�D��ױ8C��Iۈ����-1�]�Yñ{�Mn��o�ZZڧ{\��xBԲ�����o4|l��,�j�q�I�coO��������Z���B���d�Upq��K�o�:�0!۽v�z�빿Z(�9����w�b�XN�7">9d͛�rb�D�B�*T�K�x�������8N���{شY
����G�n�F��ҎO`.噞8�����_^�`j�:S��\^��y������ F�ݮ�mw�C�D�=�ӗ�����^+]0�	���������l,���2ɵEZ�P�gB�6Tv$��(�NQ@� ���pF���y�%�]�s|.����-�d�*��za} Rj筵C�lrH��n�[j�����%�&[�q�qѫQ*�� ����OT0�B{elV�[ph�j�߿~�D�mrH�����$�i�g���6�� U%&�.h�x�c;^*\�V�&vii@ �!��$�G���%��gY�Yb�A�D�l�D�L�!v{�z'tS:Y@�ݾz0]f7��"U�}=�c#V�4����Y~�>8��r���,=�Q�Zx�
d��$���O�,UM׼,��6ʂ�T��F�%^[��J�~ӛ�҉���4إ޹i��ޯ݌����[5\s7��&�Ƀڲ4�ʔ�}�N���k0. ������&_:F0��g��.�=O�����q��R�V���a����֭n0�S6���n�=\ a6���{׫O��ֿ|��{�����jD�d�����ƪ�2������Q��F���Q9 ��qo�N�;R]hR�yQh�:�d��R�i��GC������گ[oZMA�r��:q���K�뤡��]m��i9i��0�2[���ɁH��]M�6�꼽�Q5�A��P�1k�Ȼ�˺��0nqEF�V�4��}�5�v��W���w�M^p^����dPZ�C���t:�ηeIg7]�C���t:�C���t:�C���$I�kG����F��Z� K.�c�K��5o0m���t��OG�]�s���{q�G��I�\�q��_��ː�>�v�u9+ �woK˯[��F�C�q;�`���L`*�f����q��>�<�Ҽ�L�{��]��;n;�d�i!Mȍ;3spf",^tE�ܘ3�bNw`�/l��V��40��}f�(-���e�9�5_5������d���^��M^�;���)��عq��	P��N�� �9�&ڵ�q��ԛ��]���:�AT���M�4��
�4c!l8���1�HF!��҈�qI��}��իg8ܗ0�;�n�C^�%����_Jp�]���I�\��u��^*yb�K�z��~7�6�ɋB�1�ڥ�r��4�>^�j<Rt�|X�p����{�z����wxy�=�-����'�?o1��Μ=9�N�O*).����VA�n���2�9|%�w����w��^��9��(�ۀRkT�D�@���Ȥ~�B4�s"�;��j"��<�r��c���6�M0�o6|7��%j�[�q�H>�N��H��(�WD#�8A.�W(v->�w{��v�vދ��>H�`7�ᮬ��znՆ�<��v΀�^٭񸄃���Qi��^���)~����Ę=w�r�vV��.l��0Ȝ̰j�C�1�ou�~�}���fQwRf�(N"!2��
L�ڪ���.%�␄w!�*�D��7�o��$V���3?u�)6~�~K2G�hI�۝�=�A�]i%���|+,i�!�9�$��&r��n�Gr�6���!-)zA����u�3�����;�_Iwfn��Nu�/h�5Sn�h�w ̤T��5h�ϜY��ng%�f�4.$
�Qoe3�
�C����Zh<��,.S�
���t:�C��yZ�t:�C���t;%�I%�HHu�|`P���\oh�0�p:��C#��s��m�L_��輫��jڴȠpi��l�kl��t:Z�T[u�dl�#����R�����VE�� ��������~��Y�+	���H��-��l:��)�\O����V�:$×Sǖˎ��3 ٯ���n��z����Xl2Nt+5J��*���t"�%,��j��z�J�ݰĩ%��:��;$�@$��q�f�HTa��NSwp�h�9w�l�$6@$IF�w`rKy�%WCi�� ���ջ����r&�)�t�ml�ܬLh�;%�H�C����#E�$�q��U����O�rBy���=���'У����۬0`����kٲ�8sX}"��{d̎�E�_u�.����{o�  84ԂP�� L�		����@:a��0H�20��e�4�/(�� ^`��	Ba���q(M��
-�� JsIhJr�UFᷧӘ$��W'ku�Q��t:�!�BI$>QN^>z�0I%�dlth�L*�]�B���NA!���l��a@����k���4�R=V�o:�D��
$,8%�C�l0�^x"�
���� P\4�L&H�w���^�Ɖ�� Qz"R���#g��B�p([{jW�p�8�G]B�����`t:�L� 3�=�9y�i�Lӄ�$�C��C��V���CQ<m�/Z�	}^{���D����F�ts�Z��J�k��ST��.��� (H�r�m�H�RAQy�lZa;���W�4ȧ�Hm��%XԌ���U�E<<�fn��<H+U�m�lWNTd��_q<���a��J��F͝Ͱ�ty��t:Q �vd���tf;����6=��t:�ʓRv*�w;�T  �RW=���D�|C�����-��;O�C<�H�C��$���4ȠP3���z�AP� �V�q�q��2(KI� �F"�����@��,H��"E1as):�$m�3���Ծn�$�0�GL^�&%�A�0TjK�N��>�g�$y7������1������Y#������a�@���s�"e�`HOAz��f���$%��L�d��ݻE�D�� �"�1�Iv���q$¦���".oG'ٶq���ϴlQdj�y��D7����q��r���ɡ���{Y��QZ{f"M�$�ws6�NH:QV��B�|,w�s�c�;y���/��OM�c�m�h��C�ݙ���}9�r���g��q�}�K/���3������t:�C��0� DH0:Ht9�C�����,'�	$C���t:��V�/aoRk��|��g��K����ux5���&�gfs6�u%��N���C��7�9��=������Ğk���XS/��a�2�8�����پ��6�o��^���=ͮm��4?��v�7Ӱ��`�B����T�m���^��S�f�Q���w�zD� ���*��As\��>�:7`�� �=��n� @�:�3�z8%恽�rC�N{�P���0W9���4�:I$��=lxV�p9���x��0 �D�ER���'1i]-��4 &��������Z�&�$CnI$陙K�k�ԓ�>+n��[t�I$��t��D�ј����9uZ���ò[D��(a�t#.*Gv�ݝ%&���;]���v��{�^d�Oh��PjM �t:�G�A'�C�pa�ht:jri,�WS<%�C��V�阌Ս��n�M��$(\�w�I$����Ē�:<ǅ�a�P����4:��݂��a��u�t*  Z�"��D��ۢ!�ـل�耡 t:��6��N���_��b;�_�~C��	jI��;�$������@�k�ø:K�r����P8�Γ��'��{���o[D�	����|�]��PJ+|۷�d��HA��$��P(��E-,0�	$�o�
���8H�[�L��$�7u�@_��s�f~�C��e.�v*�A jj�� t:I%(�tȠ�:  ��֒��a|έ�ǀ��+��Q�lF � !wI�����I�I@f�p�H�o�l�I]��q.�C�]g[]�Hv��C���t:�C��mV�-�C���q�[k�j��  -I-i �I%0�f��H����$��C���t:��C�NCa���P�t:�7ifn�o�Э$���toM�����C���B٘����$C���0�t0�m�ʋ5$�b���$��HH~�ǁ�a{�aB'9̝&�I"�y^Cܝt�_��h���9�k��V��퓛+�l�_$�J�]�������	]ܐH�M
�I9�]z����\H8�C�����~�]m�[��PL�:���ko���/�NQu��r
�]����t::�"�}�f#�sy㛙���B!G^_7-��� t:���K�H:�������w7���wwP4&�Ѱ����n� ti�@�p:�C�ԒIC���u��z�^�jI�^�W����z���N�D���t:���a���A�I�C��-�I-�GyШ�:�C���t:�E�:9��y ��I4n���	w�����ퟖi=�<�ZԞ��]:N~��Nf�����1Z�m���8���[�ė6Tl����<�|��5����閄*���l�C$��j�&�|e�s�;e��Ցɷ�Ȭ]\�8姻yW,�P#	�w~�a�;N��UO�U�oC�3�n��rmo�}�'��:�U>�ˁYD�0\�<h���m�d 7�MR.���W��.���<DKz�L�²��䖳�E|H��%��E]��p�x�Ǧ_r�T�i3u����,��;O��yA���j�X�/���]�ZL/{�����_E�k|�v�<b�&W,�so�V|Nf���*�b,��r���׏��^r'����@?Y��B(V��]:YvL�NTB�	F=�L�@�l�"��ڄ
���4\`F�/,����q����
2zbڴ�b��s8G,��|�b;G\�_u��=��!�S�b����=��mŵ&��jOy�Nh�>���<0i��=޹Br�V����v�2�B��$D�q���������a��]=ێ�oa�W(;�ڽ��.�o.����~t�vr>��T�n ?���}���ބ }ϯ�G�Ԑ$�,�@������~_?v�������C�$�	����O��O��G�_��?����O��?�=��9����6f{(�\3���u�v'�sH��S�w!�v�w�W`|#�g\�^�!1��p�oX7�����i(����c�VCͶ�kۄї5&�ع�����]W�^�=V�wE��^�j��F�*-���6��O��Y��V�����xB	��W��_{WwW�y��g��۟;P���!���d�a��ڔS{�i/��'>�}��#^߹V�ֵ���L�Y~�: S$��d��"��'voQ���M-i�p�#��b�.Cf)U\�Э5���@|>v���7�s�aG|�i�9���V��TuRI&/#�u~|kE��Ȏww�� �!���3��3[�{���+}1-�t^�&o]��I�M<@'9�;�ԗt�9�W꽐�>�bv0}��oKO����A}wyMWdy_��ݟ}�.�x��L�݉�i���������@M��}��;+�og�~�Υh�k���!+��p�~ih�~�/+,�FD���<qMi׻\��KW�wĄ$�Q"FRH3*����oW������:z�i����'XI�5����������	��E�f���C.tV��/�YѹA��j�Л����"�]..s\)�1*{�fs�S����RS9~ ��x��?>#WBW0���چM�!7	4��-$}��9W��I�QV��j66�M�Ỳ`9�oG���O��UW=��+���a�{.� � �!%FIw]�3��uΕz�f={�9�����d����MɌ8s���x7�iǨIƺ:�����򪙉��HˑB5H�?jG/	Ml�`l��Ǝ���ոk�|s����xr��e���잟fC�U�[9��ˢ}"�h��2�+F��ɩ�Uc��l��|�[����n����H����:7H�����G���ch��MLY�F�S�ͰA�e��}�p��o׻�[�49�ʐ�2���5nDL]\�W�&/-�W���D��$���9���y��㷀Q�k:��>��M�Ǣ`���ғ�5�^|>�#�Hux�ښ��7T���Bc	'�HcI��:ty]��%����>����cL����5��&��9c`������!�����z��ffSS��^�']i��#.Y��+*>أtC�JO�E�~ʼ�hLt��^�3���&|���8'��kȮ ]|�>���at��O��h�c~1�(#_R�8�mRr�ֲ��`���:�6/���`IU����F�Њ���$�	�Dw����yvB�A�W|�UBMv���&��^ծ�����ʈ�|���E�ذ�.d�CjD�u�Pď����ک���R7#Z���3cظ�/9\`��
~�դ&�f�%Ԩ-��	͝O�K4�G��6���h�S�>L����[��� 6��~��+��C�]=���Pa����o�$�@|q���_*����f�}�ݐ�" �&{�HM��e^S%��������;��ou	6�����s{��c�_�ڢ��HB��)�y&$h��sz�o7^�Y�NY�t5�u�5���~$	i$�z��Z�QSl¥'T
�P��玲�7tV��u������e>��� }�F��m��߻̵=����fV���T�'R"����I �F�5TfB�m��e�T�'q$����8����ڳ�q��CqėЩ���P��r1eU��}��H��7g�D�� ���^Dj��ċ*�v����P�����+;�B����8�"v��u��8��w�����mT�Z���Ъ-;�u;�M&�j�L���O!!���{�{ܠ�s�]����5�����5�,�����n�9�!�  �h���lp�ȅ�cCȩ��y|e�����U����U�b빝6? �s+nf�!�Q	�kU�z��5'	9��wnk=�̻4kբ@�5 ˺��m�;�Hy�j�k��1����p��w�W�n�{y/�K1��g9�Rn��V5܀>�ئD��B�D�:���'�q��U磓�]dM�&�x��� C��ب�W9�\�w2��t�|>b���67	������'� f��tz�چbz�+�5��s�`�7�u������k�=��wB��){{މ�*�)ۨC[��G#�p��w4N���}O�U��2w7Я}s|���Ԝ���6�ﮝWϷ)�0߷�VRUR�S�5u�޻]�$�@�vf{O�)��N�o��j�/r���w.��F��묩��7�������"�u�Y��/����!��������>q*�f������	��P�;�O�FAg����,��{n��/:���x���UV���$� ��s~��}�w��
o�����J���[�Wh�y��[{��+����X�́���$�� ��y��Iܟc��*�J�����UQ*��¨��X((��TTR,b�E���� EE������HH"���� ���A�#�#�       ��C�����C����"��**�            > � 
UTVDUUB      � ��" ���X"�PQb�UUG�@ @     !   B     B      ���   A}�B     B     B  >@   �   �   �   �   !@   �   � �A�B ?
d*Ad� ����� A��@  ! ��  B  @  �   �   �  �  @      �   �   �   � �  �   �   �   � � �   �AG�    \����       D}�  ��             DG��D|             DD|G�  ! @ !   }A~�4����,"�Y' �B���<�� �n�<�������;���c�8�8888�<���<��o �8�;�1���{wޟ��I��V�B��]s@UT�Gk ڤ'UG'�ڤ鎚՛��
Qgn�h�/}�~O��z߳3(.fr��z��\�o{��/8�9��PzOw����i�3, �z�w���9�9 s� �Zփ��i��2���[ȋ�C��;�ɾ`�.�9�wQ���i�Z����$KT4L��dGf�>���#V���|��kcD�r�%ם�Y�tKo��޾� ��V���z��.`���_#Hd͝�:�����C�<hpݓn����/�G���{�z�[�s�*��m���S�~�o~��0��|�}�~;;r��J�i�U�\�1�E�WR��y�7�D�k�*л�*jB�5���қ*�Nv������6���Ӷ���r�k5�Rݶ5ٚe؉��:0ӧ���cu]��Ԣ՚��/�[�UTw1�j��K��˼���[�^�����*�3��~~?)��7�3��<�0nh�$2��Z"�����m2�1C�|�in�K��>�!�T��8 ���8*^\B���@ �7��F!B�M �֩͹��O,b��gk$�����|[��&32$bcM�Ң���dsu�?| � H��M?��	w�.��PUQ'�,a=�RI�yʽf�Z�f�d2�Κ��^�@����u 4�y#�ѕy�|��*&�٫W�"�$=��7���C��o�cw�|sx�|��M(�'�4�-�qbT�Md�uV�1c���%+�������&+T�M�[z�ee�ذ��a,a�q@�+��`Zy����73F�����t�U˧b�F��VwW
�o��C�����=�����I&Hsi���k4It�ލ5UV�ݜ �pZ�/�]���ݨ#,vL���	%WY2n,�8`�-2fq�uG|sgo����7M�;Ղ~���wq =�[���D��n.k
��%ɜ��H��/c���c	1d��BO��̺�꓆
h帬�w�lܱk�ss�n�oS�����o_�Z�?wu�6x��0�n1��<�gZ������~���R��,L�yN��$2T��U���U)+��Z�a��Xd�I;���3����dp���Ŗy�B�J�[SXW��@>pI*�^{�lPS�@	�����fg&�ٍE�fV������k�qh��Sx��W��� ���P��
ŃU��6�����y=8q��5�ĩ_��p��N��=��N"s<���tW��f�`9�i�*F���\�10���3��Pd�u�\����\;"7��ژ=s�2�2[pQ�gc��jŢ�Q�&%��Q��I��)�)�wo����޶��O�Cj2��,��P-�Na�5��7N "�L���x>����Z���d�麺9�.O��:�J27�W���]����!���}�VbԔF@_�5*�0�Q�Vo�5�Ƈ��B������v޶��y��Us�	F��,��y�laG	�V�"q;��̃u"m 䑁w����=ZM�m��T���pߵ��|j�da�3(L�ȧ���f"���UFV`�s�GF��`���ڳ�5��d��c���g��T d�UQf-�;��!5{�3L�HڔQ)���j#X-7��yb�I�Y�;p	6�4���ֽz��=^�����޻�}�U�x 	�_ߙ9�n>��SI�l³��7�n\�w���q8�y�G����O-������[��ccH��d8m����Ž=({��}���ܾ�R℀�:}b䜨��*A.Fӎ��-�ݞo~��iᯝ��wC�V*(_̮��X�8��	58���0�<;�+$��y��F�����#'�{�FI�+�U�F�����ڏ���Q��X�$ͪ��MPJD&J�g1�d�5���.쑝�8��ݸt��gRm�1���W��<�;B^`]" e��w �Vk�_ȆE�μ?�NM���ikS*J�j[��̿W��|[��ףq���]�{X����n����g�ُ�Nd~�;��)K����Y���.BA����Dsf�|t��`n,�iDG�Q��pL�d��/R�$�YT��p�����5qFj���ީ=QSս�C�5"�B�P�i�D�܍4D�������sa���u�ڸƽ0X9�*Rs��͟�QRHƃ��D�I����qq%��y�&_Т[B��biH�ªL|�4������ty���ʖHy��ޘ�0\Fr����Ȳ�kpa��+�yỹ���l���O�=����U���{"f�~��\���7*�����ߟ�?}?W�ۏ�u�t�V�Y�֮ٻ(Z�Ii^g`��O5�.e�ﲷ����	!�O����M�j2�^BōK �H� ٦�:o���l�q��ܓ[^�y����e�h�� /a�w���z�l	Ⱦ��C����v��bVŧ���O����X�LED�)QM��3i�0����>�vx}|gz������;��&����ݟ��eS*Μ��ݑG���v�S�"�S��d���6�����#xMLP(8'/I=� �Ҩ%	"��!v�}������ຽ�t~���ݬ�W[Q���v+�ߝ����J�D��;i���{b�X�z.wr��}0�e������X��e�b��nL��O�17�E"�XAJ�4�d�����>3�҉*J]���� #�y�U���T���Qj#绎�Z�ݾ���xo\��]��VŇ �.�� <���^�W�[�'��_�����%T92$��q��Q�a����ٲe�{�r����N����&S�JM7L�TE >������!�'r�H�sW_}��2����e2�P-Ö'��������Q�X�|]"�R����i�)G���O�}��d�MJ�*�K��c��1���|?F޽n�(�`ڊ?|�[b��ڃ�`�)ɾ�s6> ��_wHfk㺵ˉBC�X����L�]��}\�������~��<�e�X�E�p),�a�qQ�TI�3Q�v��T��cR�3bi�U�vi����l�D++GgTV��{wDI辢�@Q��bf�|ԇ]��O=��-d͋�3P��8b9햏 *DLȢ&�+r�Z�8�^V���2��M+M?�nAR$Q�o.d�;T���[�z��N꓇�gx����,㧶d�I���p�ǭ�K�ȏ�[�;y��)��;'��iZ�1�`ݙ!u�l�ܭ�T�ݗ�d�.3ξfr����ɼu�@G��´n��!��H%�Ѷ�mۜ��Hj����e���ř���-nfC*��(�����MTCdQ���z��c��r�$�A�UI�n�:�Փ�Wߗ�������I1��w.�9�i�x��A�w�o����z������+�V�5���jx^�P�v�>\ĬՁ5Rc7������0�Ξ%���o.�ӟw�߮�U(kT�󡦠K�՚�*&d?U��J�KYf�zD���WW5Ef�DQMD�/���F�L�b��{Bdc&2	�%J�a�ȍ��,��)i��G�TJW)̨�6ssk�f�+�^d��G��8-"�B�P�a�D�̍3{� 6m�0n)�+٨�Q�l�0j!��9kO�}S$���7�z�"H���
��́�T���:� |*�n���H�w�X��"��]ww"�^��i��3!Qj�^J@$��E�[U7?_��{��w�Ŏn�������^��獵n��vfe�@��q����~��w��w�[�Yh�T�Y�=�"
TL��;��T���΋4��)��9��Wm*V]��8IDôb�j�m[�/����oXdD�e�O�ZW�����A-���ݎBqT���]����ɪ��fa���o&ď�Fğ��<�84h�d�3
a�RC�����| �3���²�⏬N���]eov+�8C�PK�jl�Kk�܂���G�T�	��vP��)2�I�;��M��n�(���"���HFor���μ��t�+(ay��NR��D�纨���E�����֍;�[�*���}�b-e-ɨ����E�n`u96��\�FK��>���Q"C��^T� �f��ؽ�YW=r�<帤޾ �4���q�ڀ'�M�5����X�����hЙ.�����h"?W����^~��a�vՀK$$���y����<����F=�2R���=7@ۼ�Q�M'
L�̗R��������AW�'�!�yW�kE�	�#i�����ɒ��G�����GA[�5L@�Pt����'�Y��/�w�N~�;�D�۟~����~�ߞ����&v�;�I��xG��3y��{Y��]�&�u��	�zB�̸�7y#���2/b��À��SBf��g��<��S�O{����~fn�9�P0UCr��Q!��h�U�� ?���:�b*D�:~���� �k6�`~�&0��z��t�ly��Ϸ�MN��}�����7N����Y�M�ՇL��qڵT[\���tl#H>�n��=��3���niĠQ�و-)�D$2ؒ/�p��s!M�y��Y�םo�U�QL�~6g���58�3�w9|w�S�ЦOkY��m�j|q��o���X�;o�q1 	4@���Д��Q�2���~�W�b@$�s�X7�}���E��Z&�����ѳJ4ů���/e��|�yd�����+I����&H����YT��8d�$}��h9��1�J����:���;����{�&����U�7������0B��!L�J���υU�N}�Tlp�޽Ѷ��Z���DU��{�����|����{��6`a���M�D%$�� ��=��5�����&l��͙i��a�\	�E���!�$�tE8��"Z���H��%���{:ڎ��a+�%�v�մ,᮴u-�+sX�j3�E�z��-�|���Í {�n@>  ?�I�?6U��V�    J� [h{�wz�x6l� �[i� /um ffP��ޭfƷϗ������т%��Qd�t��H��n<w���)Xw����í�v������}}������Sܳ���TԢK��qX^�S��������"#-����>���{���wN�D������1��K�ذ��Q���\��iۂrم�i���gpY�4�ܾi��B�]��q$Ý������t�rQ��6�<p a��ӄ{N�#A����Uά����m����c���7�ufk��8%u��8m����&�ό����"�eż��Ypt��)c��Ξ����<�������8���]��ԮK-�e��C���8��+�#/]���9�
v��s�G��;�F�,]���!�'tnuњ�V�yx*���6��rEb�tn��.���-m�q�{e4x/>�z�޽DE��8�]��ld]�4�|�pZŰ�]!ar��&0�jv���v"�0��b�{�m�*P"qiM
��c�f,RTn�O0<�`F�u��$ږs{؟N�:����5�����?�Ws��	<F|M�Y�����IӼb�W+�p2��%�%脮���HK��I�j�Y��zv�'�����Y��%Zg
�����H����fUD�����]�/הks|��x��ַ@X��w˝�/uTҧ���ߖ���ڬK @����x�[v�=51�q�Gl��3j��&F$2)�$Xfb^����4 $Y	 �Z���s=�x���/�{SٗVo�b�+�@�2OZʮb�)ծ��<��C���+���P���l3�|g�E��v�wW3D<�z�����@�J@w��!�6��>z��v�*��*�V���S�$�h����'��~G�?��x6���~4^Ր��`W��꿙��m�����A���u!L&��x\�4 yBXs�35�7���+�e�q�0���������� QO!���W���I����A���m��3��5yuzU}vk�^[�IX�����v9��BN6�'Ą� g�>0�u$���)��$��{��0	L�!
H���q>�'���{��l�-2 ���v�n������� XV�V��u����I��0�y!����w�Ϟ����"�l!I�I|�'Xm!�
@�O�v�NUu���;SM��7\��@R-��^j|a����y�VQ
IH�����<���%0<��uP������7'@`1 �7�6��d��a�|���@)������YZ�IL�5���i�:�S���}��0�@u�@m�ۣ����j|B�

)�����2K�����{��g�)*�����3�k�:qw�ƶj�k��E�\�w����y�VL�����A6
��3LQ�/^����{����}������v�]k���n�������lV�s��1�1���`�i3��X 4�ʍf^e���/F���!��޴�?2B�>����,_˞AM�d9��i}���j���l��E��$�m'�Wi$6�R)���w8[r����T�ct�^#�j�M��U�i��϶H,��N;a��d>�d�b�@�m�S}2� 8D�fI��|�W�'pO�o�f+�e$�1$��a�Yߕ�e�B�m������S�Rq ,!5}��y���ǲ˩&��9ۜHi(��x�/Ra�k{-�r�&�d@P�� ~z��N��{��́��'���9T|~0���h�8���)��<ϻ�d��oܰ�
`Wߛ��^�6�[����Y�LN&�3̐�$�׻����!N�L�8��H}=����B�(���ouݔ_�$���v�O��@��j�WG� 3W���R Cm�I�5�}��tH��@��n�����L:��>h�����hS$��̹���v�C�ϛ��md	��C����� f{������I[�Z��t-�� ���a�<�>V������ R}����!έ��oޙ$Y�ۯ�Pc2�*�qm�� ���1>$���R0���@�ט�)%���2bM2R/���QsD���}�'�D(���+]�7�Wj�2^���yWyKv�5��4�j�s�37ҌI\�H�@p2�,�Q�R�ŧ���ѝ�gÆv�⸹��mȖ7Sˋ-�u�㔞�۽��6�]Jѩ$���5�JN,�e��l�3/<�D8�a1���W�����V�����!I�3u�>��C�
IO"�L���LKHnx����^jM�U�ʫ�N�;gR�>^�>��Ϟ��>.���d9�`)�!�w�=���H,���۴��{�=��)~��ѳn��e9�'.���%�L5��2M�"�|�I�W�H,�y���a
x��}�\a>�@�0�!Zk�N�Ѵ�<���ę��W���6���B��{��'�E��E�@��a�J@�v����PEHv��i�G��������Iߕ�<�!W����U��1��w��ff�["������8�v�U�A���>e&��a{�&	2u�a�� FU�e��vϖ�^N�-�z����6�"�a�k��ebC�R������@�>��9\)n�ۖ��QFfg$sz�é��|`S!�V��L�R�a��a�T"��8����ʏ���[���-�-�����'��$�{��[WZ�
����:!��T�ai>��������}��w�L��� �l�L������Y��x{�*�|ԆƮ�<9̑����k����<ڥ0�3�/�1�ٶB�z��8�E���<�5����߻�'~�5�nھ[͊M]j��i����a�>#�}r �� Ri�~��O3i�/�;Ϛ��Ґ:�S\d8��$����2Q������{h�nL�F���$�+{��{ܓ��>���� Di*K�
��L�$�j� �E�H�Y��ΨT�$UJ��y!a�ϼ����m���ǳy�,��F
N �� �C��W��$�C7'M�@�O��x*�7��Z�>>��\o����AkФ��?I2ƺs˦�C��]�bh)_gk���a��!���ƅLm�[`�R,�B�[Rm/�0��H��������~�H�;{u�n���Ks�y�M9���|�'d�W����f�u2����܃���,��w޾�vB
@�BU���ے_eH+	I���V_�K���.2���C���ֶtwH(��Wt�wrm���@0�^������l�I5�2�ߨ&�h0��Ϝ��q�J{��o���l��U^�9�wR�� _���p��f��ݕ�}�֨O�`ݑR��������<pM!}uW��r����,�-�b�(o��n؆A���H��NT�a$!�p�.	E�
�3ąH#��;�O�,�@��3(s��T���^J�lg��Y�54ӦD�(v���G��	�:G1DJB5�7W� �!`a�n��j"=��#P�@����o_���9y�w� qF�%�*XR��ܰF�+2GH�DUt���"J�i��(U_&"i�ɼ��'X�q�^-PǄD��>����wz��@�~�[B�zk`��Є̤�F�cª6��M���y��\`��7�끋��k������Gq���x�R��������F�����{���J䒭����N�eT��������>��/�^��=�	ؙ�n
"���h0竣.��ݒ��#6m��1����ս�J0��u�8�`�C�|�^����Is�`ٴ�켟��	c�釖y"�B�R�9�N��L=�"ڢ�|lE�L&�v�Q^�N��T�a�Æ~�{��w�p	�ȷ�[Q��X!n�
hD�#M/��G��&���y��z�;n���{�M0A	3�-�@g�W�n����|��BX���R-����!�K�SS���#9�������I`P�K�@�C�L�HZ�4;�ڏwT� e�R�hT��&\#"���F�F�L22t��}��}����!�աt�͊Af�ǘ��z�;�U1Fd:@ӏfe�>X7�͙�P�b�LBB5�ż{��#�W�j,�1��3B����0��=�v����������.���������M�4><�a*�P��`�W�tȄ�}����qT^�A aQ��*�oF�깘��T7C�mVW>�L�I��/61�`f�'��;_|����^�,^��.p��R������F���W:6�4�GGk��g߲~����y��nM�_~��e�ɛC�jK�Ce�K�^�YJ
N�9��9���������� �ڼtU0n2�f��%6��[J�k���z��E�%����
P�Cs�,c�.�믻� Mhq�C�칕v\ZQJ��L=��"Ң�|��m���+�`|,j�#�l[\gn`��؄^Ј�J�dD*��oW�	�R������on1��P�=;�����=ᓒ)��/�:_#B�
���h"/�m>?�����\[�Ϭ���~�B
�T�NN �oy:��0lΙP��冺��Z�I8�W�,�Di]O�'*K��φ�c�9�(dl��.�Dc\o��{�����)
��c�*�|͊�UDME!�6x���"4�B,"$��a�_ڮ���A 
#�����UTMU��XJ����ɾo���}{�gy|�;�)�!&���і�K����߽�X�^��G��$#,R��.��N3j��P�������wB*f�B"�hR@��m�̄�+UW�^�F��Y �F�~�����@ݑ�_�|�U
��UB6/ /���~���H|�#	=G���7}�V�^2�>{���6P�N��>��@�# %�ª���c��J	F\�"�f��m~��pfuuD�;�r���M�7�^]�bYy� }$�F@�>_�Ah)B����<�����Kl+?�ܓ�X�3Hw0$In[ns���|~��0��/��"�QD;�/��+�z.;� }?ӅG�)���%��ɶDN�u*���A��ٯ���|ԀtB�˽�v��s�o��tW�{�ɑ��{G�}��Ef�C5���!'Q�}aJ|�N�¥f\�}�ɧ��,�x�<]����[�pQ��27{���i���� 䳇�i�� �f��7 ��� ���7�>B����tV��8�!�LD�t��Jm|>�� qY�ѬS	ݚ2��hu���Y�� ~ϐ �\r?�n�]n�8���p&� ���z��x���b�;�����׫�\vwa	�=��r��@��Gb����m1kَ��s��[.���N
�!�	���d��6HC�X�]@DpB\��*5_�t�|>��;��BHP�;Д*��U=��
�}`D��ݟ�M4Iu���7v��@�Grb�������a˂b(@�)D�s0,3����A�����0+B��ܶ1,>tXЩ��p��BܷJ��*B��G��3��ȩ�Gd��� �X�̋~��RF�A@ X�o{��A�R E��۳��i�m�+3�X���]�f�ك�Ԯ2,̉�ʭ���jp�9��a���X�����_[��|���§��Z�f��c� ��\��m�kpl�=	����sr���mA����[mSuk]����k\�
���]$��*���������8�ҁp����隊�>�H"�CvjT�5�h�Q�k�b�jȹ���n6���m���}��ג� ��@�2.Y��!�K�U]��;�����G�����"����^�Dg:0'ZaR��e��2=��'����~hv���}M���)�b"E)c�k��5�����  ��������&
��E�[}�o���Ϥ��! � ē�~	���g�b��
4��>��.��^�1����f	87�5x0�Ŋ�8�1��f�7sBa:�v�|�$d�a$�0(5f��9ۈ�
K�W0�F�r����r>���Q5v$BB���x�A�����B\����'�����)�Gsb({$B���a�jR�:��盿���,v��^��$^��Qd�3� ���@�M|>���
B�DƏ�
��z�8~�A" #DdP"R�A0�(�R�1EY"� �"$�Rl��҂Ĩ��"1��B���dY�(�H����]9�7y�kW��>�I�ՇWݻ��37���u�1�L�,c�e�"��I��w���U�;�yR���Q�b�c�(8�����W��׷��>v�"o�"���\L_���I�e� �,�c��	��N���!��C��A��;X�g��m4X�˭�1b8��B^��yʕ�։��Xye1�^����]��q�����l���R'3��!�::�TN3�0�{nm����nR�4AM܅���Dy�=ʛ�|�;+����ݚ4�sO5�;�[i�h`�z�eδ>Qwו���I�e�f�i�'I��(B�۝�z���$��{34a�-%A���!�M%���VW̚�{���N����7�W2q19�Sn�W��i�o���Q��Pn����<yHC����. h��P>
�.��t^����LC�!�Z8��2�U�[3�Î���:w��]1�\��D���("1�i
H�6� �A�D�2 �,���A��}�w���c�Ub� ڪ����\[UuUmA;jѪ���G�Pz�zL�+�"jY�v:5g���]���_��������39@ {޵��@���.�s3=G��m���̠{փ���k�sr �9� ���h&�˩w��r�Ϭ���6����}�ۇ����A�b\u���߷���۟������rs�`ھ����{E�N�G�WI~�B��7�W�/,HՋd5�[��z� ʰ��ɪq���� f������<����~�vpBW��p�ƚ�fm�7j��J�����:˭Q��f�J.�LN�raDD&��f�3S
H������V��[+Ƚ�k�.VG#]kju��e�%;	=�uu����Mv�[�W.�O��t0#��^�\��9s.�֗v2��BFԄ	�γ�V�s��ku�����2�"l
s�ҶG��Q�k�:���U���v1]�h�Z��F!�QY��".�pDU�閂h��঱95N)�K���v(�\Y2�1	�Owf�v�O����.�ZY^v�Q��	�i����}�F�IƠٳ輱fo�"c^��bb�QX����j���2�*��4� aI`�����$˲���2��E՚���r���z��GN̅z�!y�1�ɛa�� 2��СAn�$��v�ſ�h'�*�Ɉ��*�)d_��Q@ ��w39C"�c6�����w���z���^񼏔��ާ��p�ݚ=˴����I5�k՘r���ww�2W� b��g�pŬ����;���¡&�ף\g�bi��4�m��D�V/E(�6�D[�۷l�]��ku���a�ba��7%tￇ���=?��z�w��6 ��dƙ��FT���m���� ~�� �B��2=�`)Q˦�C�mf��	���c?�/v?|>��B^�/�c�v��g��˚�l����Ve�������{��� �~(�Hg���$J��##��z������?����)7t&d��"� �B�\�X����2���W�ܻ��C��#�E���e�1T#J]2E���7/o���~0=�0��2��Ӵ$C���y���N�;}Q%nW&R�
AE�n9c���P�
�;�4�.3UH�gЬ�2Xj8D��%	��Nj��"!���N��X��L��إ
���K$����H��a2�"���d~��\-1�Ĥ#Z#�GD��0��s�%��B*j�(8�٪��}�>���F�%vH3.R�XK)��v�`��|�b�@��)	�~�|~ %����L��陝��L����OWu��]�Ƿ���o��;�;$�[h��k|؂#����(Xv��F"k�uH�������%�B)!����f�VԈ��OF�����Ps2*�0A"�i�T䫒��nBP%Hp\��P=������'2�q�1�����R�j�}lb_��gv���
�`t�^���pb�Ytd+2��w)�4���&�-V�]uY���2��]޻�ÿ_m�$^T	��X��uܠB8��m�BH��|>���,����3�&e�߿P���B� ��\vi�Z�����J�����������(c���h#��!U*u��"�����|����3�W30�JA�)�p����oՖ>6���8��Hm�bbE)cZ���0P��$�������m�'�1�_�������{)����a��	/_3V߳\�RK����$iʫ�����! �I�B9��{��J��T��0I<��	z���ՊP�U5*��=�O���� ��!8.p�'�R���LJB:Ž0<3v�> �  h�kJ��~�
���.�IHY[0	��ɿЋ��Ԡ��II�q�3��eK�ʿ��A$�>��-}�����@�D�d�����	EP�U1FXȍ�pg�2r
`�� R��{o8�l
�o�$�-��P�����{�
4 ����rTD���'%L�"��kT��:t�� G܂B��^�i(^�7�c������}� �a�H�q�u2�J����xȴ��/��ܸ |>w���4�쎏1mt�@�x�PchK�	�H��(���|��C�j$�@���>����|,��J�/�"�'�<N9�ICi�;i֪�8�ۚ+�Jk�{���|�>pn5L��+Ě.I0�����5.)�j��NTR6
�'4��q<r���25�Ɨ�ql�إ�?�>��E��ٻG6�Î�Y�gdϚ۶2��9�;��N
(B�A�u���Oɒ@�����#Ђ�w�C����!���Fu@�:�#)�(�DV���zG��7��l�k*�.�>� �D��'|�#��T$B��'6���j'~�ޝ����۽��cIvϕ9�)�4-�ק�j�Cwf���O�~�u�5��$��0F=ca$��-����y�V*�S�EU%�h��;�>{�>�x$�@��`J+�r�Lm1	�a�ZG�-��o?k��8He՘�sh�3z�*���uG)��s�DF�e�/lv���򚦥-]��d"+��'TU��f᛽>����}!!ni@�m|z\@?j�=�l�ַ�nBA�k��{�k�k�APD�ЁX�3�Q6����y�ۮ3=�^�����ўَ� ���C2AJkM�a^4ŇL=���n]Q=�<G�|��TLx}��?~n�ê������>���T��f��_^5�Lȳ�c�7s=;��{�{>G�������;���V�֚z�kjyܚ����Ռ/}��~/�����A�/���u"1��U�DA`��K\h5��4a�q�IIDa=�t	�[�9���j�U��ջ��&d:ߵ��e�:y���[u��Cp��&�p Z݀�e;�)c{�\�L�m�4��=/���ꚥN��E�5n
��s(|7�Ӟ�p���1� !-"�z�
̭L�N��Cn9c��e�>���B�(t@�e��Ho�Twf4�� L���%PO��I�B�&A��u	�^�E�V�#=A̷�z*k�Y��1��{���>�~{�t}ɊxG�c�%�q]b��m9�<�=�Ӂ&�'��2M
�!!�#wz��G))�/XP�i�U��|�����j"h�ΨE ��T՞��q
�� "|(�Ɗ`��4;��ϦDi�~�}�b�߿Oj!�)]z�Ȗ����lK�+m��j@C���s|�5�� ~�/�EH@�Ev1©�|>�}~�����Q�>r
0%9������ٶ�6��H>�8u���J�q�?\�K
��Xt�ޥ��qf˚H/�;����Z���C=�r	�dc�<#޺����|����@�q-��Bj(VL�
 �&��l���P e_d^���_o��;���NSJ_�<��>�O�;+.X�9��H��G�l��=��[��׿~��Υ�ջM��nb2��"-I�	�L*V�̠F!c�&=��go��%!M�6�J�֚NÑB"E)cZ���}�;׽����P��ʔ���S�t�@�7�}bnB�j�(P��r����	�R�"�7z*�V24� � �$�X	�=��I� ��������}���D��C�mӻ�-P.��O'F&��,�h0>�L��EQVa�W1�� u���b�9�r��CN/�;�m�D���Q�����}�b�e��B#D����)[j��F���M��P/N�%Bf�.�V0m	}J�h�R;y��ôqȺ��Ól��T> �ڼ5��͍1E	���tTD��[���QS�,g:�h�����p��Q4$gL�F��&�C���� �!X�w~�5&}�Щ��q"�Bܺ�T�JAQ��D|'�3����[��������"�R�6��k�����.���߾�~ ��
Y_�.�.E?C�d0x�y� A	A���ܻ�{ѣK5^����7"�sz:�MNj\\+���ߨ}���h@��0��2����a[��A�~P�D�/�&O<����n��wϓ�1mpS�;5a1�K%�� ��K���wcn7fgfU�UT���paA1mL	T�EU��G������}��PZ,�\
���9ܗmL<�cm'i�rg�v�g�Yj8�Z��^��}z���tFڋl��A{���ׯ}���lp���B ����7��'��vo���w[U�*hyȘ�T�&E(c���b�(l�D0�G��K����	3 ����<��v��	$��P5���y�7T��ص;s�+�b�\��	G�>���EO�:���7�A:T��A�T��,9���}�V�<��pd����A���;�nِR����� >��'o}|(�FS�T��zU�`�D����|DOu���~���"A��	UA.����-
tz�4I�Z��DϽZ:��,�A#-i��+$��`�*�ܱ"��W��߇�~�%�w�?��8�BH(B��1/�}��z7ۘ ����1�+a�/�n]R�n-#J������ԕ�*Sl�T���^���AB�05��u�D*;n5�k%u��w)�םf�G'ߒPM���U��FB�H
FD浜ߪÓ��M�q&�
����wm]|˻�nт�lCysU�R������$ҋ�Nf�4��z��P�SUnYv�)C0�e�n	��uۍ5�s��099�I�}��^���޽]~��Gp�����w�z�n�o��pS�����N�j� �$�zj,�-e�g�O������4Z
M<��׺��Ê���9v��B"���{���ﺵ0��2����
Ж��NF�����_}���USE
!�*!��R�5����)��8�����wz�I�\`�	'%��lc�U���h�R&A��f >�>�W��x�C�;PB�ż{�𞉳C���,��Dex�ȴ�д���ި���(��!�PW*[KFp��M��_����c��|�|R���J"h����Q�S���:�Yu˺���OI!*�ֵ��W5�Q��1sD��.?8�{���� ���x�DrP[�@��CeH�����v5�Q}+~��"�2��ٿ�o_]��$�(�A=�{}���k^�9�3�Uѓ�oFFQ[Xv�E�
�C(}���ut������t[y�����;�#d&�����둉aUɌ�e^{}������'�.�`�ˈF�٨���-���C9|�m�}��|��(c�G��mo�\�B8��a���3U��MGV��_| ��U,z�B��\vqܡH-����wf1#Ђ;���8U_Ir�E���DZ�P'az}p�DO�e�����z;�E������[��y��x����8ʀm	h3��L�i��9�4�vw���	�dL�j�1��QlS	q�R�"�����Ͼ$���I'�"v���9g��Ϸ˻�j��sDgV�@�=S՝��|�G�#�j��~ʑI	GS�1����L�^^��>^����#rH2��4���%������@C?E�K�%�IH@>X�,�jHw��c9&2H���ʶBRAd�>�:�BL����i�4��;K2�;���wRi�I�otN����8�U��bi�sӆ.�V�e�&�z��#1�I��F�4�I�1�dT\�XC˹�n%��&v�;�>%�����_�T�U~���ݞ���m�T��]F&���)|�X��R2�r[(�+�U��U'R!D߳1�%��Q�Sy�L�,h���H�5���Vr��S�<�ڐ�
=��4�v�Iha<���[�rLgPR�${���B�q�WS�����(�l�^g8|��n��w�4y��e��3{s{.ke�R�:A�*�zA#E��
�i8���2e��Y�hk]p�ζ��C��'�W}��a�B���|���k���z��Y+ Ք�5(�%�ѤH��y:���tK����Έ��K�<E�H'�1 DE����,��̐ZC�d�ݬNМ�YE��l0��*��f� �mxUmZ� ��k��@ �ə�w������h �m�������_ �;$� փ��f�${m [m �վ DDDDZ�]Y�[V��O\`e-"¯g�������}}z�����B0�p砷-���7s�d��	mJ����#Y��YQ���F!�"���qM_�m��-B��P�AE������߰;d1��������̗�7��%{������)�q�5)̵T�7��h���?W��W�I����|���]��]�2�lZu���h���2$V�l����њy��H$��`6늵�GX�5���nS�9ؗt˕Sc@Љ����5̆�+nʵ��E�Z.�B8#0c��<��u�MQ@�h8Ϙ�7Hq���H9:�r!����+պ�vW�"{#Ĺ8��"m�;WkE9K�w������Ã��`ή�6��-����M���t:uO�1�O[C&����&Z���F�ա��X̠�N�y�9t��z�u��,T��T�i\<b�F��De�"E�x�����Z�Z8gn�L�6��
��J&�U�#�z1cvl��w����*0mbѝXή��Aq�����`Y�}5\8NX��f�߬����	)��������o$��`��o����7BcΣ���>�'�OvEz�4����K�_�#�G��s�v�wR޾?}�����\}�����ӹD���w|��z#�P¨j��T	-���O�5�V� K`��[�/gq�I�����y۶�|�~��m^��g5ƶQ��+z������+eWL5A���W��?����sX�߽�D�j�Pn�@�,��x��.��mR3��n�kj�j�B�{�Iҍh�jJs���@�T.ŢP#��zu0ȑv}��U)"LU]y�@?Ͼ���_���׃ SƉ9� ~Ն�K���^��/���3�5SE@�O��rJe��P������\V6�»znJ�d�HU(���`�	���Z�
ABkm��a�E�
�{g/D-ˊSQ ���2z�R���������ۚ����/O1MID:^�ݶ	�\~����vX�}�|@�3ߘ��W�\�[	mIqQp� �A|wvi�l}��)Q��`3s�%
C��ܮ�Wo���߁� ~��MdA��*�q������0�ZS2���+�{ }d�Ǡ-BZ�r��=�U��h���j�G/,���\��'�^/�/G1L�bKEJ���EH ���B��5U�ř������?*��'~!1�Rcs(�]����у{c�g��h a$���*ۣjbR�0� �"�H��yX�%�qn���{;��nyV��r�#�d�&�\�����M�t���g9��]Q�<��&��c����7�u~�߃n��߾��� Ôa+?�  Ȉ#'r�����s�S�n��?�MD,;�:W�P%���������;�l��e�z�w��~$�ty�|��,�Q�����Ϸ]jaIC�	�&��n��`�>�.�T7 ��4_��蘃��9!�*����G�����)[*�rꡖ�qlx�DZ+6	U_#*�����*`tM{�0~>5ȓ�����/�:(H���S��77��U�B�A��!)�bE[��y��yi���^f��F`X�����1,>vXЩ����n]R�MŤj�C��߽#�m�,bRQ��3;.�"%��7�}=ջ��P�`�٧�@��wB-�I�5�l�	:��� �M���(���/m͘�y�:9�}�~{�}?}��?�������ÙGW�|���I	�H�@f��m�6��tE" �)"O0��Vc$�y'�s �RJ�($Y`
ywwu��Hp�&�:b:m�bYr�lՈ��S�ܛ�h`���n�3͍��fi�i��9��G.(���:�(�ڎW�,q~���������#e�?l&P @)J�0���ra�� I����n�5��/�	ƘT�+�`�XL@�ru;�:����l;���F��	���c�]�s����� ��sI��*PDq�] ��D�5����/���(WP�5"$�)x�<z8T������~������a��C	k�lc2#:����D�=��p���p~���������A�KZ��~�>�QR�d��D��fKU�bȈ큜��(A5 ��ͨ�����,�iDq
B/��}��D`���� ]��4��6�%�3�����1I@��b
'�?}!(�����Ӱ���Zn7�" �{������|>�C>5��)��~�A]&�[�ۖ���~�V|�,$���6����5!FR1�n��A%!^�n��}��孶�+3��.dp���A_J��Æ���萀�)��A+ΜP!�y_i�;���ȓ����t|7ٝ���}�I,���c*LU~�b��'�1��(��/?|��;�~պ�לb��,���t���С�����=�Wy��x�_��$�N�VO�����W1B͛��{���9
6&E�{e��a� {D����LO�c�I��*!�H$�0AF������$=��:Z��}��������k�=�t/�bF ��9jaة\z;��?-yD�5�}5�X��_�0o�m~�n�\�!di�s{��c�q��=P��3�,�X�'�X�[�� ba7��s��Q������H�~�z����������� ��uf�Y;(�t��T�3��Ꜽ��uǨx��$#w۫1�hA����<ˉ|`�:�h�%��u�nD9J%�rǆGw���T8�=k�w�#i���Y��˽�����8����U&I˶��b��g�!@���h�9��"̴F֪�`s�k��`k�ؓ���F�"��-����{������k%����G��T��D՛,Q	��:��k�Ͼ��n�r̦,���D�ZB&e>R��s�K�|dY8��ZKɊ?I
�ލ�=?}��~ ���yHlB�dȸC�G="l�/%�?}=�כ�@���Yt@��"/'ɕ2��_�{>|��	!��{ܟ]'������~��(ԇ�P��"g�ݺ?�Wy�|�qP�lf�f�
�p�6�.k�[�I<����ݼ(�D%.�♅%jm��-��L_}|�|E���S-����	���� �i�7=kQ�����/%xl��s����-���^�5���Ɏ����ln�
D����u|k+�ޏ����5b��#1
���15�o=5�����w�w���nqXi�ɋ���y����h�ē�$�kDW#I߃h�E{`�?_�Bfk"}��&�
Q�#�N����&7`_&Cũ��K�fl��߱�P}Ǉ�2*�#n_Ջ����oh~Vz/c�`��7|ś=\���m�����뀫����DHR�d#�M�� m�������Ѧ�/WR��E��3��4N*d��׮H�<�z�ѳԄ���Nn���E��c�ND���/��g�����[V�2RQ}�R{�%��
	J!GН���C5i.2,�'�u�̢�� =������E|�}Њ�IPa���mT۩��ĚP����FU�F�f�W�J��L]5sو$0��	6`lr�*vjo�;͹\`q�	 ��`�3f^�]ЩD��_0orn_o;����g�66�ی���Q�P���zD�Zc%�$�g�F�u{*�8�Y*<��Aj�,���t��{�gwW^e"�8XB!�/KXj��L?���uə4�\�E��g&����Gm�隦��F��Sh�w4�Q����<3/���EG�Z�<z[5Y{��� � U]͍՞J�;�͐��r!��m��}/i�ٗId \vŹe۔���앲�����饞�,ُs)�Y�)�I����Ns	��ƽ�Jg�d�w��2~GOf� �2���}Z��sLj:���������_��]�s�@<0�>���ԋeWϞ�n��[��&� $X
AER}w������|ֹ��2���i�~�����g���=����u�S(i`��V��E5���|t�V7��F�8ͽ�Z�,�3�L�I�Ti�/6�B�v��|>���y��7S?I欏1���{�J	2.P����Pfu��\\sDI���a��q�S3p9��<�-52�Ñr��oG�| ]U�&3hT�O��:)�$��T� ��P���s�B���`C�x��>Y�l�Q�����SԆ|��^��@1_F���oKkS�uke�U���O��$e��Mă��&*�4$����6�OnP� է|��{6R���ر�4��,���P.��;F�{�x}X���@쟅� i�E����������n�f:� }Mx��6���y���޼�󴝞V�@��A���8���f�X�H-��An�D�5 �󛋵�)z9�2~^�7��[sm������5{P���K`���SshDWfȒ(�p��a^dԥ�u ����ť	h(;y�ua���鵷�z���t	�Q�(Ґ�I��(�#"fS&4�7�t�F�8"�Z=;ױ�Ϩ�:��?��,#T�"f2.P�ж�+4X�J�ĲD���@�E�����z�}���EM�x�J��`Y�/oꏴ�SY�\�n���銰�P�:>7����0	�̀g=����x�-�,�	�$�+HQ�� H�'��ʠ|�t�8�i�@��,���CH��;����*�u��G/l�z�!4�3	ߦ�-�I�H�+&T��S�A�t��K��z[�����|׸��������ήZ�#'��dzс�:s�t9T�eW;�z����
��M�ǔ�n�Ƥ�s��ߗ���9��w��;�� ���n��d�!ۻ��wߗ�]�w��N"�`�#��UW6Dv��?���>{�l�S�p��v�s��~L�P�C�>��̑ �l�(�g�-t��b��PeGगG�3iQ�Д҅�m�q?|I�����E��WOG��{���^��4��4R
kK��9�m�G-RYc�� ʓ��frE�97���k��O�}���I=
+��W;�lP��=�H���x�9�����?�w�9�饗��|ő���S�'�M*tS��{{�| ��1��D�pD�b1~��N������Ǆ��{0���"R2�@�CB�Bq-^�φ�`�r�����p��5a��Br������"O�w!�"ȕ��X̓L�P���@�Г�'�E>0�	E�Ϸ��|�:�� ?<�3��7�=S�Bɾ߁?Er��YIg}�/�h���F��yܺd��RD�$Dt�� ��`jk��?^�B�f���w;6?��ˑ{�<ϣ$�`]hD��{�tu�$!2�������[�o8�K��ޡ���Ek4Ĳc5`��3LÕ��:h��Rx9��{��.����ssV��0���2�:j-��]YPc:]���1n�fW\�<R�¡�����<���&KH+Jç��Xj�+�뭫e���b#6�آ�<��!��K�U��#�lt�SԷ�ៃ������ffV� {ֻ�h��/�����$��n�lffR�$��{օ�\�w�s� ��ց3�����Ud�b\�6�"C��v*戡	:�9w���R�?��vB1����ĉ��!��#Ӝ��.��j��+Q;s'�V����ܰXח�z����с����,���DPѹ�FV{v����Or�Ώ.[:���2�&�׻�-���Z�G�d�W�Y��nc�ʐ��c'j�
膢
P&����C�(Z6ܣY����u��)7WUsj�g��Q.qcn�qX�4�S�:�M��v��4��*ӎg�W���X�/�Ӭ�E�CYF�9*���V���#WpݖԜuֳN����&�n��I���������"��r���Y�vv��`(-�6�i�\���Vm`��Ј8M����,x�St�I�occP;��5�����˽-����5������$9������t����l�Hr��*KZ�*i��JB��05�ߜ~�w=���SĹ����>�����I��F�r/�)����({�}��뽷u�5���̝i}�ZL���{\����r��$	9���nn���B��Q��J;Z���"ɥ�*h�Z*w1���J�]��?BB[������s5r���I̸�b� V�8[
I�x�
��\�ҿ=�o�}������W�v���������8�e��#u���;:�q���o1lۮv�-����`'�~��O��{����xQw�����<'O/=�f#U�n����pB"��&�n�G�d�+r�ӏ²�£B%�d����Y͋�&�\�E�=��k޹����4:pM!'�bB�W�X��=� ��T�8ꤺy7"���PF��DGt����k��{�l���Ӳ��.BFFܱ��|2�ݝ�|>ܩ��+ˍ��|�ُ�Z�}��}���l<c�~�E���TTЖv壝,Q���&��v�]�ހ�H��4��p[D&�� ���qD�99����Le&�-�ÈS3�L�0$IrT�(�S���8"y_/JBڈ�̛�}Y۳�Թ�ӬY��钜��	:�GO���*����O�����HJ
@F�����9��I�
J�� ����U���E	�?{3����%'�&��ù��p������+o/\��fŤI)h��S��� ���6'��Q�Z�B�q1�~����;��Ї0�s�P�I����>�bt�1����w����i������b��7)B3-DO��\O�x�޸���U�:D;��Ѓ�5�oX�\�F�騡5""$2(�7��Ps/����j7��LΪ��O(�������A�7!
�iz10$]��MĂz�E��l39n��HjSQG`�"3=<���5a���D
��1JHb�zr\�h@˷�zv=~��P�/��|���w�>�y�g�E_gv��F�A7��T�C�r���(���}�h+0@��*��kwxOl%bi,5՞�	��a���'6���U��ߵ�ִ�P�Q�)�d�.�m.��L �)"Tm炉tr���.��O#Z[�s �����|'}޻ꨳ$Q��O�;8��׻���W�2�w{�DO�	�5R��:~�΁8Wފ�k�Xm3��2��X���-��.����/��r�v&(�$#����ıR��
����<�!�����&X��C�"l�92�~�ow]gU�"���b#9�jRq?A���ި/��g0� ��LA+�q¡xCޫ���1�_�6���3 �DY����u�:��G=���F������Zr6�Uʹ=n���vp��@�PFG2DXb��#��? t�>��˦T���:(z}á8Nqр��rU����H뉭{������i$��$�y773=� ����%|���Sj�6�Ѹ�8�-�JB!�˰��dAv�	��q#�"��Cf��e
����{Ss��UÑ���<4���y�wfo����H��K,����
<�}�]DĐ�g
����de��quS�O�ќ`�{y��d�CM2���!�@�K�������=����z����H捧2��}��Q�O}"I�D$��ҁ�Jt��h��d�^����y��zc�7#����=Ii�%k�m�KrhE�>����U2�7�Nyޮ�cޟo��&,��#�SJ�������}Va���������Ɵ����W�{h=�����طP�*�L�D�7��Y��n����LfI�V�R�NR�����}�{��]�&�������������ͯ.?�#��^�fجq�A�]�������\��A=�c�RbO��j�(H6��$��!�,�0[P�6�n�������>������>�4��>�gd=��{����;��NU҄뵻<�q�C��Y8��n4k��߶�����9Th����[m9���$"`�IXJ@���'���6w`s@f�pN�a_�uP��R8��X�f�S�����ˠ��΁�5�U�f��-����71�1��77���v )5-�2�$d]����E�i��E|&�n���b�}F��(`�P��M$�x]ﺄ{��4��Fv@de�{lp	����Wc��M&�-�ÈS3;1RhD����z;������p�hUP�wT�#�1��Xdު"o]��SA�{�d���+�TXKiǷ�g�Ae}��T�6~w�t���p���c�=苭�߸��Q���{ɧ�\��(a���".�|?li��ѽ7yUUU�W{J	2B��9-���Ϻc�kz����t���'}P�w��^k��>��X�sdI5�І����F�=�ZJ&Z�*ި���q�#ӕ^��|��0����O�p�U��dyO{�ڷ�U�[@fZpN��҅��7��\E&�����Oܩ�
��Du��ȇT�"k/&h.쑨�)���(�oy���ܨ���1A]��C.Z��K�b:|�ߚlm���LR��?�5�!����C?A���;�m_p�����Q@�!�&�T�T�ۖ�F��ս�+�v���w�'=o��t}�����RqҨ-̰f=Q*�DE{�F�iU�a��~���#���cXd%T�UDG��M�Q�V�_x}��F����$4lޘ�8U+�Oj̪Qb@��׹�o����ZD�;ŽLY{z"'��Ҋ.bY�뚫�;���WՐ�!z��Dş�#���Fk���f��j���p���4��eaT	5�Qd��]���ئ�2�M4�%BE���{|ȳ��Da����"/��ƽ	��׬<�g���`��.�T}�IvF�M~-�����L��,�2�M��5L�$Q�3�ݛ׽�xM8'��,�X�.�l��7�`���`��y�1U�	"=�|���l���c�����/�،RC�zunS�R���vGw���qHz׌���ݸ����&��PG����(���O���dƴ*���3Q�h�t���;�@��%[}wov���.6���)Jܩ�*
�3BMA;-c3��:c'&�t��ӵ�i�;�N�g���jۂ�KDv�[c9���˼���3=���,�!
�� �� �,���ܿv�EX��)E�P�N\�z5�2G��U�0!��C0.�Vvκ������ϯ��^���'6���荤�쒵��7'�yWa�!�Ad����nO�$Q�Y���l
ՆM���~���BR���4��\�5SJ*"TA���l	Q�L�xTB�IȘ�������dvn��DIBTi{�H�+NL�G��ٛ�o�l�<�s�[LfI�W(R�A�P+����{Y����~�s!��l^�;6}ƥ(6r׼D/
gTɥ&A"���;���&J�
�͛4�����l�6�!0Ip�N�o��RC�l��i_KG�����c_�:�y磿7���n��T��DO��A����NLOyZ�{rueع�	w7�c�fr���O����t�n�����Bћ��1؜t��X^����������v���ly����0TUm����	�y�Xd<��@L�RdĻ2���/���U������ i}n�A�ǥ2&\����^s�}Z���3�]s�O�Fn1�����ck�>��{xhr�Y��L�bD7JR͖(������'�y;��[�au!��Է[f!ҙ����
���R���B����DM���Q��+s��wq�.dr�������v�	Ҿ��|~!�lD��PO�"[֜�HCh&��zs�F�c&0�$i�������~�z��h�{��ct��v�A�(i�^�'Rœ-'�9�}��R(i1���7(m�r�Q2���F1oO@��_�z~��d�򩙛��L�+(�O�F[��r�4f7�r�� ��|�QL�0YBd���Rw����v���"'�1x���5}�`�¬7U!ArE=���6ۂu{�ۻۂ.�"��[�h�"����H�SL�QnG�&{��4W��U�#Ô� ����|�f�lV��L�6�ǡ�&fZFݿ�<��w����w���<�>��7��k�,?�!�QJ;ݬ�x��ۏ��y�����Ez&��Ul'ۼ7��Z'�M�U�`���J]��?s]��F^?Dw��g���ji4�3a���Ƹ��3�3�D����b�&�޽�1�vv���DD�0Y�J(��:~�́=jo�W���O{�� �ID��m{�g�����a9~�Ȥ�J�|�0�Cw��_��>2{K���?��H���k��S� J��|��M@�LIN��2�b�-���\�����wF�S������{��yoi��Ɖ^y2���իe��%/
?_A�؎��]����=v�y3O��_�;ٛ8G�5���[ϝͦ�����)��#n]�{+�U���a�}���[��sG>Rh���J?S� �������Z�eie}4���L�&':N�]0�
sWu��.����N3�9ڞ��vn�w�,���{�E�y�C�*��Ği����Ė����=�#��~����ޥi��?D6�;@m�4���҅04Ρē�N%k�~3�i���4�N2S+TCeV�ϔ̨md�a-�J��(��,r�{^VJe�V""<։�"݈�[=��������#���r�BDJ�\D4��ۚ""&Bz��� �M�o!���f�6��s�<l�ކ������~)-�;�f{����h �m���������6m���m�g9� ^�@�@ ��̵ <  ���cw���͚��G*&�[xyW2$�B �80�;	����l�݌v�0Ae�PXMB��4({3S��T��B��"aB.�2�\dS�I9��L��J(P�:63UT�\�^���:Z�q��q�CX^�P5���.{����q�Ax��� �⛯f�eŶw�9�m�i�JK!�B	0��s�<:Я h#4DD���n�X�I�7a��Z���v�+��[k���	�j]�$vs�gM�9�e�F�hksɹe�ɱ���=gi�C�!������Nq�z��NdWĲ<���<�N9��u��N�Kv���x��D�1�l5	g5N����Q�]��7�V���xfv��q.�Cv<�p��NhշN��r��sv�Ԧx��7h�3��DO:�m1�f7]�C,rp����.�ŵ�xt��s�e��sI�f��� ��"p�z�����(�!��W��`Ƌz۝�q��l]�{8ɽ�<u�x�f��;�6��_������A;��ܣU6j^8���"u�s��PJ ņ1�'{ɂ����_}��q��ǽ�|s�-�.�S�{��q���~�C{�u_����@�{��TQ�`K����k���t�y�������{ġ���JQ�|��Մ{/�s��$q�,�6p���HkP�FKZ�(`���T�Z�� � �5�s�uŮ�����p���Vέ�tS�ѝ�J�_7Z���a	%��������{�ʽ�}�ޑ� ��v�J��kD�~���H�?F9���ћ�����n.��n7T�b�fEB��^��S�N��͑'�[|x�m��ĺ;R�F��\��O�`Q�[�Q���ʪ��^TMc��E�u�D0ˀa��a��&�1z�؃gr:Cz!+6�ڎY�}n�h���P�LL?F��W<F�pN�Ej�V^M;%z-��i���-9�EU�D���\d��v�m����T@�Ƿ&=�����;Ƒ��?�)�p����G9i��G���.��_Y��6��#�ҚJ� �󪋼�G���:g����19�ޞ��}�@���aH��$�<w�u��m���	�H������Z�o�/*����n0����$�}�����}� �I����@�Vwt�����d�TS����r��Sv�d%Yv�s-�nexv]��=�yj8��Nh�G��s�ӺBV� 4e�meMճ�_���c�$'�YqE"ōV��s�{�؇RVrIZ\��n�\� H�]��#�DM0��ۙK��0�Z�l�	4�	^�j�&�i���1di9�8�J)x\��HD��tZl�L8��"\q�7}l���8"�Y>��zj���~�!�p���5�5Y��dT!��i����\��h�?Y���d����m��2ʥ
[H7*Rû�a�F�s�W��b��A6��7�4B�Q"�dғ �]��8��z��Hz��z��Ә�w̟���x��3Eӳ5"#3�/����*�N�D��	B���-.� �C�ӸFVg2��ܗ+�����=��$�H_(�iͿ~�nxa�Ei~j����v�����J�f�ٸ;��m�#==�=���j�[�\]D3Jm���[$1B-��#r�'(4y�:��7V[ye4���5g}��u��=���H�����ɔ�˪�߷]G�m�)VV� �HK��_��P(�-7��O�Gn==���G�X�(X�Q���M$H�v����z}U�'��]�22�ɽ����Ng�7�����a�R�:"k��B[p/���ތ�QO���b��,�����s#U4�M͟|���10+�}A��+�	�س�z�r��{U�ľ�)v�%�I�P�����X}�ݱ�
�ϧ���߭���qlݲ��[�������Z�s�[LfP��অP�7�1�aI�������\wg�qE��;��� �����;I�80���&��B"��X{���}� @���M����T9#�m 3��JK$#�y߷_q	����������]��"��p�j��-.�D��ߴ����L����IvKe�ܪ�.�Mċ��ʋS"���RFqRG�ǽ`ޙ��@����e��C.L̴��c�q���ʚ�Ƽ��OC?Asu��{۾�md��(�~"4&�%)���h��d����eh�����:���f�,��#�g=�x�����M!����M�
&X�%�m�FY���3~}w�������z;������fN?| ����t]K�^�b�>��4�((Ҁ�Ɵ�s�x}�ݽ&�q�KI��Y�H����f��-#32�SbEJp��9Aa����Q W�p�l���|�cݺ6sa�f�,��h�����L�헑1b��&@��8�%� �H�$���v���b�!�b��X�ŭ�r[�������M׳x�޸@�U��`M�b�!����6o���Z�%f�	T "(�=����y�$�YE�޽z,`����;r0g��������L�7!�Iz1��Y��`��tC�¨\�L�1�Ke7$����N�Dg��Aҟ�5a���t��~��]��b��0ܦȖ�F[FO�WmTN�㝵�q��־���ex^U�oh�oi��"\)&I����X�'�|{P;{�AL�;j��[He,{$�!�q&nd�����+R�B�J���'r�Ӛ�@����? Df�8�;���:/Mz��B��E��a㣷fan�&��>���kn7fgfU�UT��m4��Ta��������4���ON�i������Z��$n���46tt�la�]�Zs/j��Y�W��F6U���s��=����mr���wc^Y.�*�uʪW�iOa�.F�IR��3����A}�} ��	P����LMq&a�ܽ^�'"b��F�><��*��vϢ��Ժ�aL�O���_��	�:�Ӑ���Ld�������� �����3N���ɦWCRS!)���ިʍ��^���]0��8��'�
� y�Z����:r�L@C�xt�d����^4=�R�I\c'�}�S��J3F)�T)Nv�wo	���H�2������|O���m
�\��h^>�J�		r��]J�r��Pm,y��V�0�E���C�؆�8���?A������v�y��y�׭��Up���H!P7t�*A��9��U=�'7R�A����y�{����l۵\�U�s`���iG�_�tD#W�-���]k��󯞾{������y�.�����)����*Y��qs��w�oW��k<�"��E��a�����NA0�� ̏3�-�b����)�b���8����3��RzyJ�aB���ND�H�]�exV�u-T@�\d��!9縺y�}����p��Q%̎��TY��{v�TAj�������NǣO�Gv9:��gJ[��R�12*�W7�^��xe�'�>���EU�睛�1y[pܯ�e� ���z=�в�}bgR�

�b\DFA�}*�z�n���%�0kS����5�˃^M���Q#	���@Pl"0��~>(�m�:�r���B�Rķ���,�̈́�H�J�NB!��0����ښU�$P�$(�!���$w{w��ff��m��PO�hm�%s�uޚ�Ved��(�?&�~�TX-����'����������v��~3����
�e��ə���wo���4o�M��2<';z��T�5��=�b�vრ�M�)�3�g{����d�g!gc��roU�����wcoH�[:�lB����DU�JG�����M?j�)��YEY�Z,�X�)���\���XD޽ų�,��7���^�P����X9BH8��5!8HY��6�TA�pE��c�=�e���E����՚��Q	)�1"�7�P=�Dz���gDs�O�+V�B��ng�����^o�L')2*���@����#c���>��L+�R
|�Rp������omE���H(��Ց'M���߯W�;�����������e�u�@.�g�[ۋ����D�7A�W�!�0��p%P����w�h�V��8F[pN�El�E�ͯMۊl�u/zNG���ڑ$Gv��PG��K�-�Gsj*���D!��N-��	D0���"�*1s��?oc�Rd�b��0ܤṍ��\DM���m�R1e�����ʁF�q��~�8��G�����1�P.���Dȇ
I�tܕѬx| ���\~�U~bH��VGF�>���n��ȔU鹙�r��C���(���N�Q�w`i�ڴ��ُz��4��c���R�L�T�#�5W@}��@�
�¢����b�������{U�>,�7�"!!�DB�
Fd�L�FDWm��U�DNL�J蒭�ۼpv����:�h�T,o��}��=z���[mq�Ls��k^Ec����y����㌕��ť2R�J�W���bvz��c|����$���~(�1���"r�o�hb�j\���"�7ӱ��:�/ҁ�0K�ͺ握BG\4�� 4`A.֯}g���B�=n�1���|̖���	�I)*e"Q0jP��"�r��@���5�h��g�����A���E8Y&���"��/�m�i���>PFƴE��9��w����r<�����_Q�݁~RFt�G�[�_@<�MT|O��ێL��XZva�*d$$m����{}�B��x�g�O�GZӽo������CE�x�Y�JDÁ�>���[��׿R^Y�z�4n�V��B-�ne��b��&�Yi;�z�_�++7���B�P�0Y'�$V.I�����0����@��H�� �Bd��ёC�w�>)��'}@Pq�����&�0�ݠi�6���R̇�I��&�^H���H{z���yx�{W!�M&!�{Iw�ѕy����~�d�o36�usy75��1��p�.|M�:�CL:βN��'C�wA8ì�,��R|Bu��F�e=юŨ^��~ʇ#U�q��u�D���7^�����TO4���M �Z�kI��B���(�6M�]AB:��U_n&U�p4W�e�5I��h�!g�{b8�y�C>9��m�L��y[��/��4i��8�oڱ`�A�RZ�|H5�k���Fq'�B�Ϛ��c�{`�u����U��$�o�9�|�9D�#F+"�X,�}�@%C���$ zN��|���EU�f6�V�D�k\���Uj�ڀ�]6�U	�9��kr�j|6iv{r��g7/Ͽ���o��@�̭ =�Z�m���s�Ns�Ns3=rI 2[~��ʲI=��{և���$�s�� {޵��������<`��
��_����vו!ݤﻼo$��Y��
H(N�4��0IEC(g�~ϳ۬�V���xS��EF8].���oLy�)o�]�2�Ÿ 4��R����c{LDAO����:.OF�ӳ�L!���pz�9��#�7�w������7a��6z���'O���}�~���̝6=z����(�{�-�f��C�1��+����h�v�QW �k�0�G4�er��%Σ/e۝�vh����p;B�R�����̓�������]/�Vl4sێ{wo7S@9�Mأlf�="ۊݕN8�ǅÌQ�>b����^1�J\�����j�W��`�ј��P�* �����N���{������F�C+W���&��Ҷ����D\��#j�&�>�x�g���.cb�6��&��}6hā��̥��=�Z{��:t+Jgiwx�O1���˓&Ҽ��~�5@��
j`LIi�yB)�U���M�=}��c�:��Ù��K��۽����9���W@׀��碞%	�4�T�b'bf�"D��Yz�� zj�ŽEɊ�í����\*u | ��>�z����}�}����0n��;��I�����}l݃f���O;Sg�r�U��^������|��jESd���^g�`C��"�ӜW��W��|��e���&��iHH-$.$J�q��3�&,cZh�R?�	X�a�?%[�a�g������В�y��A՚c�.dm&JQT���X�����Y�#�G�#}�N��2/o�2d�2*P�;;m#����7��N����,�\������$D�NA�G���������]�F������3Q�o�!=��&����DQ���GH�w�ݑR�{$h�F�\�0�,�!8��A<���h�;E_KG��k�q#�|�Uّ.���$3�l����ʛQ�����H�zP�v�l�x��ܑg�^�%��Y>~���n�W�y˛���G�D5�X��R�}k��?T=��fx�S���)m�؞�^E{�����j�@�Wy�&�R>�H�!r�f�ϕ���G�#3޷���b��>��������n��d3p��b���P�܁諾V�v��^VFWz���ݝ�4�P<�����>��~U��Y��O�{�>�Ｊww��ƐkFl6)�� ��s�����\*�	��w��AFQ?�(�PW��#5i1�~�7�ݠ��Ď����ɱ����f�F�Z��=!��z�������+�?tz���Dn7������2�`(S"�a�u@���{c ࢢ�'���D�/���1�*d*f
�N%S0D����6ۂuO��}~@|>R���*�> tJ�V�؂�q�vu�4n>緯���!w`�~Ż��D�	?F�غ��V�T�G6~�6�����
*�������w��@�L�q��Vgr��|�f���zdI�nFD��#.��zh�.>�^[$G�ԧb�v�n�.9��n����~�=H^���s<�Q@���4a���r����&�\��POz���Q��Z�ݬIz���`�J�+��Kv%�9��s��]@s��?{� |�e}+��q����{�}Lx8����������F��w5����P������{9��7~�2��V�5T��2*��螪��(.66_�~�y�	|J�o�]�  ��k�˲Pܜt�օ�q�	�g�cW{;�I<�"3*�n��(�0Z��� ɖH�ڛ�Wl3	�ʜ�pЈhAk�a��i�bl�%�譎�rsծغ�W�g6gI���Z�76.�<S��9�\�.Up�Gj�$� �������_�c�����0�D�KN�T ~�b���=�}��޽~����W��HY����栋��؀&�18���z�`�"�|U#��g���P� "�L�Kp��4�էy3�R��6��
�ʡ�/\�~�Gܼ��SF�t�_��s��[ۄm�d@�f/�>'��+6c�=w{уc�񨙏��		r��ځG9i���G��z��s�{_�o5���I�S�å	�b�����Lmfh���}'�f�H� ��roU��Y��x���W��!��n�� �*����������O��cIH�j"PXE@)�� ^�j�&���{����1,<��\��L��� /��O�n>I,.��	%�ӕU�G󛽺:�a�{�=��K6���]:��Ͻ�׷׿���щչ{il5X[�[*��F9ѝ�ks;�Ɗ�~�oY�n�FS�I
.�z��=�.��Gi�a���u�~{��TA�pD�zf<=5;�ӿQ�1e�N-�&L)�(a�K���wfu�f���O����Ȣk�;���TM(r�2ې�T-=�� H��8����v�lM�l�� ϖ�;��*����������#�r��6�/xONb��4~�8�!7=*�T[q #~�<d�TB_+�q��a L&L�-�Ze2�k���������֟d�Bd�ߛ�^�j
�0qFےR�l%
8�r��7���T	7ˍ����⛊���zi nM��7M)Q&�V9ߛÒ��X(Y05vI�����1��$u�TT��^k�mHn+��F 20�]R�d ,"�HAS]�yX�!�	�?��{ӅR��x�U�~����K^���*��������sKM������߳{�m?L�e�
&\GD
��6��*?*؊8|;}^�X�EG����g�Y0=��`lTA5Pb���o�q2�l ����a1�~�9�^���Y����ܑ{2���&��f�_�]�&����}~}��zݝ� ��8V���4;��OڕЅ�\�R�B#=�&|dJ�����cR��$@�(aJ�ﶗ��@�x� M�~��S���=Kb\<������!�DW-�c�~�n����2��h�.�/%�-�DWUө{�Zr.(���	1y���#8�!}}��}I 
C�7���}�>��f;���O��~|�ϙ�f���l��r�a����F�~�{��Q�����3���?u��RY/N�)@���h{�>�r}�ݹSP8ח�d=�n��޾��g��_HX���-H�ّ����O��B���7b,.�H"5PaAA8M(,�o�5�Ef�Ŧ��SJɥ�$ΐ��>���ּ0�ɸ6�|�g��ߧ�󻙽��(���Q�dGNG����=ۘ*|ꗶ��4�Zx��2dUB�"Ng:9������+	阳��ێI>�6�hf��	S&\͘#��t���y��������0�*�%���/D�iL��K������*�����D4W�^W�[;���=�ޕba���̚�_;�������ٷDR�h;aND$E�M��=���¸�3;T|�sϫɀ���`K�������߮����}�;}�;nh9�s,�^rg��vm�܎�[c1��:7<�/TFP�n�-h:Pճ�=wϿ�;n�����@Y�+.}���z��
t��q-7NeDGc�A#���!A�?T)���	��$}��{p*0EZ�Eb��5�
�z���~�k��Xd�A�$
QD�1�I�^�~0Ft��Xb�׺nf�?O���!]����"!̄��ZvW��UD�.9�P�{1�+?Y�[j���sth�;�i�t�0��P.�/H��]�դ�ݠ��lY�:5��idj+M
&��FI��z��KKЩ�W�7;Nk��+{ܹ�1�1,8��\�؊�	�!�xh#�}x�G����ֽ"�k[��������O����Ѕ~XNÚ_I�>��է�֓2`���� ��:�ɥ�BI$!@m��@�S=������������x�4�[y�j&&�ٻYL�(I�B�W<�fʍ�g�s�k��^��G���l������{/<���O��᠊��\vk�Si���\��#d�#(-7�J~��#{�=���+�uH{iu��#�)C1�5�w��S=���0'�f��$��P|>�7�W}�'�j�U1"Y2H�+��~GH'���7^�6=�����a�̭�0�)*-D��;/�sg-�,2F���Vgr��}y��n�L�!�}�!�P�mM�Z{�;ˌ���v^��I]�:��-PE�7� K0⳸�vn�?Y�a��{������ת/k߈��(�ḷ2pcZ��BOݚ��0��X�^^;�>�G�5�ڑ�LELK�ʑ$�0|�|O���B��U�k����Xq4��;��4��64]�};����Hj�׫/gN��6�����a����;U���;���]��WuW��
a�O��Cti|}�� ����"��oc�������6��/u"�e(
%H��#�����;��R6�b�$���0Ez&��<��R2���.T eB�F�o����P$��E���S��l!�a�&#�o���� N+r�ĵ����qK]��A��p�@�n/�h�q��'���'H�N��y�bd�����-}m,С��sJu7_IY�}מ�nA�=G��1N���f�8����.���4�+$�1LD)J�->���?~W=_7vh>�,6�A�y�K��;�����٪!�R�^�x&>�e�7[��]�j�r�cb�T8�����G��?q�#N5�����Dr̾[��=`vi>-wF�[�
�C㦓|��cV��|�淮��_�cp�!��i����&�٭�u�������!�tC9un�����Z ����SN*Z���͹�m��v{��S.�j�Glj����f1�bdh�]�g"�+!&(��������\� ��L�ۊ�A�=آhT�a�T:��e1����PP:�
<�pe�ŬˠR��{3*��|>�B��!�'�B��`��YD���-T��^�9�,O�"")�
d�(�+�"��i,b`)�N�=�]v�E-�Y�Y�)hI����x���M[m|�����s�M�  ~���a(�l%m    6�  �����޻��;!�@�-�K�r@���� 9�v�Vݛ���.�����]��:or��/5�,���l������nݡ�F<�g�W:����!|R(��(��FȐԍ��j���h�E�q]�z��q[k\� DEk�w�{��~����u�׻�vn���f��t-���9�i|=���ǵ���9.O8��|�5%�j��8�V�/�87��دH=|WN�v���vp؀ݻ�â""�'DEY�+a�q�<�E۠�uDkq��[/\���t�l� 7M�4n�^wZS��ȋ昸m�1��z,�賠zLv3��ʯ4�ۥ��$x/M��[0�\�:w;h9yQнû([��������M�#�`.S�,L\�����է#e���$��87Vڝ��7P9�6����l�vZ�5��hlNjؚK<\�v\�h�Q5$fɉ�kV��k.�,m�ڴ$BRqq]r��\�V�/'6ч�V��l�r[3C�Y�D�.d�q\PDD�wx�"H�j&mC��fZљO�X7]K|C��L���^�k��[�b�`V�m���G��v�#� ={��c���N�{ �bE��}����Cfh�u�������G��{��n�I�Xh����W�+�瀄��@���!8Ž�1rǻ�}�>���7�̺`���f�5kMYF�ׂ�i7� +E:i0��L���� Qٽ�/��x"^�o9ռ���]��_a;��8��/�ww�CWX��5�3ylPm���L�4�f�.^IJ����A��wB���*��_��I�B$����v�S�5CtBAF���e�\w���g{�������y���2JI�D�����	�Q4��gquD:�t5I)��1F��Y��`��rD���ѧHde�Zl��ۻ����|7�I5�$ΐ��N��d"�<E��Y��Z���ۭ]�q�p�[�y��f��F��&��=>�di8�(��jnj�<W*�*a��OJ2!�Dմ�!�p���z\��������\s��}CN���	*\���E����W_��B�$��{`�#J��ʝv$ff�z90�DK�F�v��	�jd{�q>��t�j�&˴�9��S��[�Tӗ,�|�}���Ξ(�m�:Y��r�Ὸ�����+�o��y����\�m�U`y�ݥ]%a��6���������$K�I%M��fwp�@���m�T�M,6�"q��I�*E��x�M��&��%M�9��F5c�ϊ��͌k塐M̧����.�*�4q??�|�wP	?i��|
@D����S_@����銇L��\P����o��j���l�]�25"K(:1�"�M�^��"��Q��~�皤�]����/�U,�����3�\�XP	>.R�	�jc�8{T�:K��{»z����=�}~B��:P�0����/O��hq��sG��g�76C�Լ;�~�k�K&R4�
Z]U2�*��x�?B��������Y���瘻�#��͞̍p�TR��73Q9��h4A��z���G�ٙ�D�LaG�ÄckI�*���4�{�젴�!l:�����P���qRF)����~�WZA��/i�]a�.�����@��F�}��}�D	:��-z�nVaFU�"	����s�V�%Yu�.ܖ�@WxuL��p[,�2%��p� [?;=��V��5/�ƹCnZ�i����;�����gd�`mBF2HS2�%�B����[���Yb�K�#�Mq��G�5���h�����d��yn�1�R���,�$	���s�YۼA7p�"�Z"�RW�����)*s#���QS�P~}�ix�!qg/�;T�l�<�PdO�gv�*�ɫC�UF���	f!Q��5���:�����2n��,�����Ĩ�J4$ę�Z�g%��?zY�xw�ۄ��C�n4]O�[h��I,���L���ii�6�i4�ejF�10׀�Ef9���A����D��ā01ޡG�T�"mu{��K���o�K��J�d��;遵Q�A,�<wv�|�P`# �$��>f����(�#^����]�4�(H3wr��>'������UUVM]�IH�1y5��Wn����w׋\�d�* 
al�m�E������;�f<�_2�k�#o:�����JE�eC!D�PF��zE�Zlb�==���~�c�PG�4�)�!s)s;%�eHP*�������ɘ�'�	�A?N�r���LKv�t�����ӥT�T�&�q'H�F��h{Y�B��I7_4�(� ����##"�R]�Z�)Z+�%#��2!í�yZb�ap��J���D��^��$`;(@�f�^{��f�<A��Oĉ~>$��Q-�E��i𽞮�������_�ݑ־��΁� > �nV�@����NZnb'�`���>|�}|��I�7녀!�����G��Υ*��$G[�*ӸY�jU^���~��5�ٰ&��#WVZR@ 2���+m>6F�zM,�$Α-)s��I�G����]Pw�}?i�1;��ȏK�&�Ｊw7��ˎ�@���K���fE���F��+�M�$���]�0#%���JDGН�𳚴��4��79�Ծ�f�hn���� J��Ql�R(�S�sa�^�6��b'�[�����w؈DY[(l�&v90�DK�T������{}����\@�����Nx��=y��Q�4`$���MJ�O�;�Ǌ8E�p׹�bXB�R]Z�n�NGMIT�D[�����v�J�S�{�� j�/HG�`��/�0;�>����A�����n���pKp�Rp�������;����D	�+�U��ovp�;�����G��_=�\����U�^�v�]�n����e��	�I��y$�i[���bPqZ�8sӼ�NG%�u�Z)]�ebv]����ݾΰP�Nv��P� 	� � ��[� �8:Y4;�1-H����Z{i�9�O�X�K ���3e⚭݁�Z�����|�o���/hTF��U�è>�S]����R�H�z�d�^+A���I�����0E���Ճ�'H�^���͔��AB���D�D
�>����+�Y���NeGӚ��Q[ٜa.2��.dRq�R�!�Ÿ�#1�ݾ�gV�5n�}$c�G?V#�Jd�r檈���z+�]���6D����C#� vz{���Th��u�ܘ���
%�{� z.j�c:�Δ���)Be!�D���
D��ҏ�Em�$��^����w{���'�^��kd�(Xy�3�tl�	&��BQ5Md�׹��s���7��`j3}��$����v'��N�cp�y��Cx�:yڞ%z�6�(�r������>���߻}��V�JI/�$�@��뚶��;��C>VR�
Ϧ��d��M�F�'n�$t,���%It�&��e�2����Emm�go��i����: � �t>�5�7���T$D���(��w���|�n+����H������艻ąh*4��Z��m^f��O�I��ݳ��#qd��e��v�}q��K2W)�9ɯ��&0�4~�.�	�y�RV�N�S4Ȁ�0_�!!{�KN7�Nk�Qˈ�s���}����'{.
6��t����?w{>>�tZ��a.��U���~�#�jA?m�^��!�)J��^ꁠG�����Y3� 'ڠL�����ADa��i��yUU�3L�%e�7��1�>�3��뮝���9Tq4B��)�Rؤ4��&2e����q�U��9���ZA��o���]4�%,�L�L�1�R��=��	���|2�{��f�Œl�n�,���#�*&�5?5컻�F�q��U��0GBĆ�U��̱���V��	H�)�*��?#y�0G��&��m�)�	��="<����>�oP����a� �;>$�ztD8�ʉ��Xfy�lSm�_ms�J�Ӻx�O1&�i���#�vx�
fn����T ^����DH�Bd�tD}󥝬iG�NN�#O�������wěQ�� �3��I�@s���5�q��e]@�7���6�~}���f�CG���#�|��l�A�U�f2vB�_y�����u�߳[,R�<���YP��	��f��i=��&���hϟ���У���b
2(@�=���Dzr, ������7w�| �ʯwh�S�L�C���
CQ3
��Z�����~��}���������N���5©����Y�� ��q!?W8���N&x�rW��gr#WTv��1�I��DD������	�B?I�y�y��$�-T!Ի��#�h7J�D�'5�!�}כ��t�8�EE���YTC����ﾢw>nE��	R*��?3y�Y�_���b}� ii���o#HDM�6D̉�J.������ݿ�Ԫ<��|x��ʸg�|ϟ+��0�������I9��h��Hw�]m�ܼ�k@l�ke�z��/]41���=��{�{�3�v�-��	�S*
G�3T�=�"�2�XnIB�[`�rqN�֘�6)1n��mW%l��/A���V��b�1A.^���2�2�|�^{��V諥&%����@�� �ʜ���as�(��|�l:���L5%X0c��?w�IUf�T�=�AҙA���f	Q�7�}y�H���y7:l��tl�Y���((T�!	���	[���@6��4�.��q~���4�ӑ�;���&�X��N,;��25�%TR�!�{����C*�5����H��Go/vG��.a�!K�.�H�=�Y���,c�y���v���#
!e�a�y�m�ܗSJ>���uǏu� H��jg�&�nQ���Ut���bϰf�aԡ4�?���|*D�����{f��d��8p_�#��k�G��"�W,��� �Mu+�~��M��>o�<����ƅ%�����z���7ˆ�M V��]�SL��I�Bc*�I
a�4�C�j����]D�S���d�N(������FIͻ�WMqf�n���k>:��ӭ�HM[V3���6��d>�I�i!ש�XM2B��!�Cl
JgPP�Bާ�)���?|"%���.a-yWۀN�������9����e��څ�$c@"0BH���S�D��F�8��p9 �g% �Җ�_,�h�!�8fYH�uU �P@a�����,d��qXV>�u��{m�ya����(�|+�Z�:�N򷌚+:g8�V�)��ʾ��Ę�!�ȳʏ
���I�>O�}�?�eˤ�Y�t�:�p���غ�j��}�a�����W��.����ݻ�;�z�I�۩q���:�5�֫fݩ�uV�Z7d������3�U��J�ՅSj��z�w7������/��@�̭ =�Z�z���s����Y =$��|ffz�������{���   v�ִ�^�1�3�����Q�C۽�����s�;��x�4��fj�W�	���UK��� ��A1�HD��	�p�V�r�&wVF[n�sً�<2�ͥ4�!�wNg�M��{;k��� v��3w���{v�S��7�y/X.���s;�2*��h�����燻q=�S:4Vfl-�Ċ�sT"m�	��X�[�-5�]�ʭ[J�������mK�]��;V#Y��h{.�KJ���%5�NH��x�`�'� ��������f˶%��
*�Z�K��Ǯ�5�-�vk�\�v��eR�BL-��+̏+�@U]!,����+�.�z�,�UV�ڡ�;��=ӓ��cU�4�6�2�B#eF�]MBA�P���j�����ᘨ�Twu��{y���%������Oi��~���*x�*�&��{�F.�«��	q9��qu�I,�2��D�"���aY�0�j�و�ZU�{E/2�sCˮ�Zڵ�.��'w��ү5�5��]�w($�d3]��f����w7�杠x�f{����}�#�]�%�@���n����	�Z�!��Wn��O�V����M������ջ7 ��%�g�6�^�.� �Oא5T�2*�踆ˇ
	�)���S*�l�ۣ�mHv귷����!sG���״����z.��`n�xdك��uu�Y���ΜcEw�Z�3�ǽgl���� �Y�"��ai�.�b�w�k�v��n�/���*��~gwj8�ҟ��s�΋������ȟ��lr!���ʛB��R��>5�3��#��<l�d_v�������1ei7����&E�aI�k~�΍#	����&j�͑�Ύ�kvV�)�����#�7��AI�X~�O�<p������w��d'�q5�"7�ci�"�X�,��ؠh��I��x�}ׯH;�c�r.s�z���Eo��5��}5"N�{d:X�J{3��J�/�_5��(A@p#�B�U%�+'dew����������v�*w�P�ĥ��A$�"��tx|8������留��}W�;3Yej_��٩���hqb��}�:w�Ý�R<�[��0ʺ����
?A"
�y[��`t��"E�\��a����c�z!Bj��(3����W3²�ߵy/q�q��5��'����*���}����X2X���7!���O��H278��q0�Br�}��r���{z"���D!��LAPك
�L���GV�гg{pE��[3^
&�}2fY	,��d�b8��iJq�<d�I�c6�5��^]�.��.��2Li\��r��!�́�{�(mLl�*�}�1���T�}�ʂ�I��o6����ߟ}�ٺn���I$9P�,�C�@����A(�C��@i��\|��0>2�NT�� �D�> m�mp��"f�6�믵eu�w}�k;�U�^�vBON(����ŅT�IˡT���������{9��L��{��(��Uª��{��([�8�ӑ�=뻷y����gK�É1S�c�D��|���R���;��|�$������>����5k.Q��½�������o�=���Z%A�P���c�+Mc��z^F��3���.M�î�uP
��ʑ���Z��g����,�0�����l�4I>>�ᡢ�~=N�ם?�e�<�*��7�b(�ļq�C%��\�3Ez��f�f�mu@��7nT#��L��K`nZD�X|�c��F��MJ�!���Q	&�7oz�I;ٙɕ�UU7��f�z��zވ����߭��_~������b��d��Dn|��[�nZ��\a���`����͛�&N��� p3sǯ����]��6�L4�6Ј�I�r��1T�����7��f�G\�
�F*.$�T3�G����=����׆����9B� Wef⍗�sw'g��K�8�3�_��q@�V\G�р��RAb�N��;{qB��-������wq�3�N>PT�p��I���u�����$o����)m�dF���w2�S
T%���G#�L�C��f��J5p�*�'L�ۙBj �#�-�w{����J�F�ݖNٮ���.��!x?N���R\�v��/	��Q��ٚ@��F�&�P�8-|X������q����<�S3��݃a�g/�޷3#�|����Ȁ��(I��@�)�����(�m��	��~���h�O>~\�e�|�;��@=j*�6�OF��ˬ�X�Yy��3q��{���|��b�U���DQi���QDX���X�S�o2wZ�;��캻���X�g�=:�%��s�>����>�¸ϧ�Q�s�O��&.vGlz�zǪ*�qGٓs�]��o�=��ưL�fY�EOU|i05�U4�|��s;j����2c��r���{N�#Q	�e]�I�z�#����/�S'���G�3#�F�iOfc�Z5Pr�=#(k���&��Lfm���4�4�I��(��C-���zq�r��F»�2�"\��Y�M���I�U�c�8��I7|����|<�{a�oYmmӚ�&���ϯ���ʁr3�����5�����%Law���gA�mpjM�X���u�w����)�Q�$��ƫU7����$J("�����v��m\�U��4�8:���F��$�3�إQ�b��ڞ���� b����*��&{#ę/N�����WO=��bR��q�#���6|2�����"�<��2̴�8��a�O�H� `T��L(fd��Cpb
A�$���`޶��MN��^�f�e�(�����\k0��a�y�*î�!�͑DMl\�*�u�^����>��e��V-M�uQHЅ`�u��Ms�y��eđ��N��vr�yϡ�rә�Uk&4�w� ��">�%A\*1���f�6>ֵ�@X/����c<! ��u\a�B� �湊5���y�֝���V�y��v!e4YA��!�H����j�0�vɟ�Ut\kYbq3�C
b"TT��}^.&8��I�r�ݟq
*�_�7�vܘ�N~��;�����Fztͅ�+�߱��{n�|�����O��2�7�\�ǻ	UU>��v���)g,�P�'�e�B�۞k��06����U�:K��$�|{W)�J��6���׳������:����������}^˜���[����qa�nđ�}�0��R �n����u��ծD5F ɘ�L�}��;��cw�4�ˋ��>���w���gO�.��Ϲ0�v{�������kmʕ�Y�Qf�i_߾��� a$��6ݓn�� ����jQ/'j�݈99�	�-�*4�p�8d[�pi��[��%ؐ·�<|X����k[�1�M��*c8�X�V�$y��^��}ߺ�[Ãn���M�w�<mcxHD��'

i�i�!enX�olIj�֣3�,EE7��(R����;�O�F����c`Cݰ��$^XO������Mđ��#�=��>�%0�!�0Rb0���������P�b1��#�=��w�W�Q�nN�6�*�z�}Q��������M��G��fg��zE	�1�?K�D�ϻ�!�5�g�~�����X7f����kZϕUR�n,3��v�p��S�gKf�ڂ|�&�A7�;���Nl%
a�
g*mVϢN��]����p��P$��l�D��D�)$��=�Q�{7v��7��v�=��z7'�HT_}.��X2��~g�Pȅ���� ߼���bYr���ї7 ��T��d��o����z���܆��]=��m�vm��=�l[�v�kjw�������}�kÓ�sU��3SyK��
B��Ջ�z�/YX����*cD��P�&��E7����)���D��y�4�w��+�9S�*_��xQ�&(���mQ"�y��K~�0���r���9�����D�����H�G�>��2��m�^������O5:ؒ3�#���4���Ne�j��{���OL���|e��e���C�M�T-�)�%�\��ǻ�D�*�W��߳���޶�~�T�`fR�N��q���H��r��Ã[hb�̶��p�X�>[9޷��4�	b=�
�=����7.S՝Wy_;&]t�'��J�0��E���C�����A$A �q�~��˻������nNOn31q�۸tl]1A�_"�M3P��_C;n�wm�;z8��ѱ�{׷�V����}�UNw�	'_j��Uo`��@�&)Mʵ9�s��O�8�P׽�=��f��6��k0K�u	�+�/g3>�AʯD��[�좫2�mx�v{ۣ��y�k3�N	J$5��ƾ;H{�MS>a63�"���L"t�0�.
	�ȤO�]��Zj���n�t��±rk��Ͽw�E��{���cc��y��jf�P���Sz\G{ʶw���#dD��5H��|����*�7Q������O
q&\��y�ɩT��xdo���L9����څ"�_z}D�݁ ����x����5�}�s�s8�1=0	��)d(ɪ	F(�!����@ �u�s�������N�F+{��O�F�3����{�^Oi?I�>"H��\B#��5(�L e���̃���!H�Q��]���Gt}A:1��[�'�@|@X|f$��yʳ���:�����τ�t^��_X��2hmGI�����.M@O��~�i��8*��S��@3u��n���@	�i���Fa?Z���D�ւqT8��D�=��F��jv����BwbK�RVҁ`�y��E[�*�PS
iXR�U��=_.�\l�*X���TM�. DT�i�BV�5�����;7�\scV�e�~Y�w��GNʕ<T�$Q�5ۇ�ܚ����y��7�&TRH"S"Ȱ* $ˌ�O�r8sۑ9��e�VS��%Q��H�M�ؕ""!�i∋y��nRU""�""6�֞�{)���#h�����+&v�.dd�v��i�������v�Y�9��U���.�A�䛐 s�������{�w����Am���{�׽�>�9��vܥ��Km�ffP�Eޯ�   7���j)�j�͗�q�&��A�9�;!�n����L�	d��0Pn�SQDš���"@DF����\�9.o��&N�k����������ׯ[����DCgf��s��Y������F�Ma3�tz]�v�o5k�P ��3�	.f�t.D�G����!GL�-���(����y�������斲��k�y'D�DD@�#4mZ*�웜�aƮ��)D@	5f;wd"�pl]��@S�[6( C����i�5J,��\�+pcN�vX�Ӯ$̀�����&�݉�i��Sƹȳ*�ꮹ��K����j�a�M��f�Ƀ[,�玴Rn���ȳ�Vg8�+<�rK���˃i�gm�eM'	Z���M4��c��L)�9];��F���7h�v���v����T,��J���tjqۖF���C��9-�{f���0`"�����ƵvuE�ov����w��f�Y} ޾��{��L�^�I{3��nߜN�#v�vѶ�Z��Ye�%��	~������9ӎ�-A�y����J{2�/+ש @}��=n�����nGw�|�܍i�Y�
- Ռ�mA����w��n���v毉&�����9�{�vO_��-{�sp�<�D8�b$K�J���t�̘π��[9
C��ʀan�2�1R�]����%�=U:���f�b�)U�~�LB�a�����&�O/{���6�^[Gk�K:z�巜������Ѹظӣ,J�ɍ����j"�y���OBP�1M$���Q"B����S�ﾹ7s(�*�O`�����f��+������h٭p#x���^�����F��Bp�ʝtTZ�z�DQ�$���ş�z�W�X��q��w��X����!�s x����1�5U�=��	v�I$�л���
�qL{�M����Gk�\EO�Q��F�%�m�F`Hjr,9Ψ�z�`��?r⊬˝�{�U���~$���D5P����L����	ۋ��tz��������O\H���#3������{��}e��X��8������}���;�޾�p�|��A��#������UI�o.�Q���"{*ukn6,̉�ʪۻzQZ薪]0[IDA��L%CqY�����L?j2��L�ăͷIg\�1�,oK��;�!m�U�o���/V�����ܕ/�1�';��׿}��ۯ=�8�=��z� r������*/6�s��si�<x�k����5Pnw��P�����A�/^�O��~��j2�H�ez����y���������|�d����@ivF�1��a0�j=�QBR�����q1<\Б{����Б�Cp��zI鋹��1?F��^���y��3�SVcJ�4��q�?
&����ڪ�� ��A�n�5�Ɉ���z�ֹ�ϡ�+1kS��݄�L6D9��Sq�}��|6i�*�s�J>�ގ�f�3�=��¦8D�2b��A*jb"[��zv$�����TVn��]�H!U(D?���Q�ל��e]��ڸ�&�^cI�/@x�HuJ��Z���>k��s���E ���X/᪺/����VCE�[;�Y�,ۘ;�&n�4�l�4�J��n4a7�[�L�p�p �/b��#r��`�A=��qr-qq\��>�>���ޏ}��_�=�_�n�>?���f��q ����:uG�2*�]HM=��5r���w0	1�1�W ��&ce�I:J�if�+Ϸ���4���~���=����ggu��&�Ne���D�AڏG���y)�f{�����2��ZvU=��WR�CD�"�<2�s>��z4��$$W��uW@�-v�ؠ�z�j�TU2'绱���'��,���)�%*p�)�S��6���on�N�5X)�pry^���М/DW�rP8J���K�˝��ﶧаF�m��x E���D����O�/��'%ڝS���?|s8���S_r_ c5�531s�lw�u���[y����o����g�br����R����I5���,��$�/oo�	9\�'�Aݱ�͞��������>���X�E�9����}G<}�O�7z�D�Mڸ�FY��i����CXh��ސ>B��&�]֚�;O7|z�w�������0�X���Ti:f)�0{6�*������A@��a��hC�^-�u��eđ��U
DVk�\J|�@��z�NT|a�A����껞�v��F��xe�������`�T��P��Per��"$��ǽ=������tI$M�˔|��
7�� c��.��f������pָ� �����ʯ����n�ݱ�b q�Oe�=���N�ū c�*��E"��mYIu&ך�	�ӻ�1�s'xS�������EI���
��~���n�n� m���w�{����ࢠH3�r�D�YSjz_J��NҶ���I]ц�ZEш"B�PPA�ݪ ��ݑf��P�9�/�a:�0�ꍮ�&�RP����&"��|f�Iq�I3Y������5�ʎ&�_���B2bc]2"d���$lTnV�yJ�r6z��n}��	"զ�L�MIn��o�QB��phS���\}�Gd>:�:q�`�A̚�1U ]nt��n�c�3N�7����8\���U���y�����|����z`�٫/\=�����ޝ������G��I�k���=�$���g ��\������z>��Z5�0��v,�[O����ۦ�x�H�n�n��5ݰ�mW#� ��jV�e3��|������*{rI\)1�.�	%�^��ǽ�3�W���M�*`QQ�vz8���!������������������Rn1�ns�ץ����YR�l'�I=1w3�F��B@�[�����6���������?ov�F5��힚�	�������|�Ѫr�;z��;v���M�n2t��'��z�'{�}�}Xf�(R�$۫1蓞���O�Vv�Ir��+7��R5����p�����]�_h��&$��;���ڳ�:�s=���Q�
�$^��,;��������{��ׇ�ۍ�,i��/-^�#K����8fs�G7r7������l��|y}� J�"W�������a�a�PHfA�u5�W\��Q:6��˼	R��<�%�6+3߶�>�{�������n�%�	�1�ɬ6����c���<w�Z��6֤�A{���i'P�ս{AUQ7iޢ^�Pp#|4�8����I����/�|߽���p��:|���a�0I�C*;�¢}��7����NJ[s��3�b�4�<��K�
Us��"F'��{�]��77��Ģm�8�4��UL�|��كZ�V�WfƴkEvl�o�0�{���LOC��Ss4�����Q�e*�mMՃ�L�B�$��N�����o�qyB>�+�[3��F!���T�%n��M�-�J%�π1TuN�ŵ/:v:x9#�v��wu|O���O�Ji�hC*èΏ}t� z�-O�H�ι������˯{��}���)��\w�,bp_]�$
�N���9t�o�L�״�=�f]�(��WU��}�6=�����Z�C.��ED��h�-�tD�ʼ�ft���M/w;�dt��±rk�Z�T�TW^�}��	���$��M,P��in=Q${�?U�g���5R�Z�5&C3"��Lq���P9�	q���{�0�2�;
"J!�����0�'J��*U>��9s�2�2g�M|���D�m2�(�4&&J��}��i9n�Hܥ�f��q���q)�qf���{`w���ww��Wf��^
w�_�w�_T8�N�)�&��$�{��A�za���}�!P�O�U�D#t�=gu�Il��B�ɕBy����f���g��9��,�z�Jȥ)�x����m�ː��ͽ��r�ێ��q�W��r]5F>�+s�3_ծ\D�����7��o�|\DQ��D{��;�`u�&�o�=�&E�S��Xa�pPذ�:�����wf �˷)-�\�pS�}��㚉�ܭ�7����\�T"�		e�u����F5и|>T�]��"kb�,U�B]�Y}�'g�2r�K��L�MA�����v�O�����87�.2n$���:}���[W��I�C��H�2i��Ǵ��;��{�]ݿ ��1�zUt^�7���m���O=]޺��Lx���z�� n>	��>v�����P���Qr��[��s�b���A�M ��izSUÏ~v�{��}�HY��$��2B.��."
Q	M�B��f��̫����I"�	b@�[54��8��oG��{7߁�\�+e�����D�'��P,�wk�PV������^ch�C4����	$�PXU{1cv�gZ�qe�E&`�E8`��9�q�_�$�����F�1?F.=�i�
��2c=Zn����E�H�!�-�<:�K/V�X)�brj�'��檨�TXsiC>V�G
Q��@9�{{�L��pNۭ��ʱG���?V�BP�"I�Vc���2w,i}�������[�y�*}^ˬ���s����"%9���gbH��y�{��UPo7��y�Mb�1"�B�N{,�E]��ǻ�i����zr(��������op�{`�d�l�0S��cj�]I����9�s��A���L�67b�UKb7���N���5x��g+׻w��e��?����������?��$� ��I  |�M2I@����PB ���Q�r��$� @��
�i�@��@$��hXBI N_�XI$��!HB$ $$�
�l�54º���$��@� 2w����?��w�G����w�������>d��%���룧���^�������?�$����_���G�?��������/�(|��$� ��h?������&��7���?���I �L`H�  ���,�/�?��!u�)?X?�?�O�� ���~����~���@I$ ��������?/��~�\��q��r��>C��L�-����s��o��ֳFC��*ϟ�R~���ߺ�g�����,����I Ht� �����E��H, 1���a �
A0���D�0H �`�@@`�A ���d���H0�H !"A��0���A���! �d� $ �	� �A H0DH�H!H$H1	H,�`�A ��A ��� H1�	 �$H �D0�R�bFA$���#�A �@A �$$���� �# 1 �A��H  $`"�A� �@d"A��d` 0	#�$"$H 0	�"A��@��`0���@H$�F �H$	� @a��d#$`$`2A		$�  A�� ���`H�BH�I �@����	�H0� �FF$�A��d� �d$ �`0` �R
�A`1����0H"A!�H �H�bF ��H���@H �`�@` �`�R�ă�A��0D���
AH0����P�E�"�H��X
H#@D�$B bAH �a�D��@QR1�AETAH

AH(
*�ET#��AH# ��@A�d"�(�D"0��� ��� E�`)����E�` �E#�$��	 ��! 0$@D��@"@d� �1"@F � (@P�,�,�$H@�0��0���!J�2F@ D�Ā�`�!� �@H�H    A 2@@�0��B��I"$!B$2 �� ��@@"@@H !$�@a�2 @d� 	H��� 2 � � � �@�$  �H$��� $�H���0� d� 0�$I!# d�`�$�I�H@H� $�	"$���HHD�MI%H�$I# "H�  	 A ��0� 1 	 d`D  �	��@d� ����$`A�� P )HC# $$�!!B����"@Y"��!!�� `��`I��I! R@���B DH P��`��X� �B
HE   E�#E��$�" � Ā� � c R$ �2H� 0� ���@���H
@b@�	B(H��I"� �H,��"�@X�I�

A � ��bAD�H0		@H�dH$H1�b�	�A" �$���@B$`0`1��H �� � �0��H �`�d"A $� �Ȁ$�A @d�B$D�"H�@	� �d	H(
"A	�A�	�$$ �H1 �� �H1`1 ���	`0H �� �$# 0H�HD�$� �d	D��0H"AH(�A������}��������̿��o�(�$� .���s��,4�܇�o������?��¯����3����������ӡ�_�!$� 4T??�Q������>O����+�6_�%L��B�_�0[������:?�M����G���~�?�����=-k����������~�I �Ь����W�a�����G� ����g����I  ~�$� ������|�����O�sp  s�3އ�]�J/�w�?���  ���Bh?���s�W���c��J�FeP(�T��?Xn3%�ʁ������O����҉��\	$� ��?�⦿�?����>l����I  ~����7����0��~�P0��'�?��/����
�������[������?���������/��9�
)�*�$� +�?�/�=?��?W����S��|C�O@�H ��x�������A�g��4x`�ϧfW�1���]��Y���l�7���������>��=�	ݞ?Ȫ�G���W����?$� ����v���
�������g�u�>�(�Q�5�����}�U����g�~���C��  �?hx�1s�?�ɭ��k�������I$��O���z,�^ݙ�)�K�������?y���e'�9�����'�O��C��C�e5��=��H�]� �r	 r}���ž�
UT�Z�P�I�%^E��]�#�P�ѣ{K
 ��i	$)U�5(�T)�AU �KQ�_         I�[ZZ�i�4�*�ʕJ�UQ6��١
��D֩���QPYZ��V*�m��c"R���Hi}�z���eJIRP&ͦ* ���h4*Q$R�T�Z�*(�J��J�ARѵ�RJ������zb�� ��T����z�w�i{i,�^����k���^����tw�u�s�h�hw�v�;�Nn��ٕ����#M1T�S�Ҕ�)JSާ��J�)%^�'yJR��Iy�� �1� .+� :�8 t� ;u&� �. �rjkf2��#vɪ��Q)  �p ���  g��x <������磠(��� st� ��@n��@	�4��F�j�s���UB��R� �9�PQ۵��AzN��:׼ 7�0 �wj�;.�P�ڜ ;�^��=x]�%Z���8�)՘�U P���z�tӲ��M	��[ ]m�����(wS�  t%۽<a����i�ֵ_ ��*��P�@ϛ�H��o8 <��� ;q 7T�t�'P�W8�F�e�]̷ pց�WmZ��l^֕@�j H�� ��2���� \��o��ݯn .�o^ z������]GAk���ޣ�z ;zmi����8�RR  ��}M����t('8:Ѻ�; rC� �W;��m9J`` �� 6Ir֍D��] ��튢�
T�G\ ��@�N�:J�p mف��^x��x <��x /��� 9�޽@ �,զ����1����� EEQ� \8���8` n�N4 ӆ� pp�������8 -־� ��z�@�                 �?@d�*���L5O��JU@   USm��M=UT��i��`5< RT�� !�&�MREMmF�A��S@SeJ��� �������y��Br!8 ��A� �2���6�0'�`l�o���Ѷ�08��L�l��*�m�`t������l�0�a��˗����?�y�>�����8�Ce����b�jE1��j�A!���mon	�T]�	�(��/����W<nVý��f�lt\�k��vY�y�M�sF���fF~�� ��������ܐ�V�e��]WܵV�������TR�a�s�����;��h:FĆ���޺[�x�y�{��fM�,ŵ����]N�m�"�@����AB0V[)���X}ʬ�%'������wq�S���:���g5��"�F��4���p+B�K���Qi�`���mD�d◪^K#b�����]>zJw���j�r��pCF�,ø~ՌLq\�ák�a)��%hʱqX'c:�n
c���Һz�{lj��T������:�����n$�mC�iU̺5,��H�y���d�hiH�*B%)M����GhӚ&��{{q[Z�V�dn��!�
��0U+.j[T�ӈa�3EjF�($��;)���r�fba�T
f��!�j��u���u#-TwRi�s������3�܊�ۦ��n�������92�e�ʷ�W��wd��Z.z���vmy�ql�f꽏H�sjJٗA�����l2ZE ����m�EB���9�,7�v(�/m�V/pZobw�mY�*��T�I�F��I�m
�[,q�hǓ+�9��.ƿ��R�jwn�)�$���D\���v��ds�US�.6uVb}4[[SМ��<�K��m	���l�Ű������z�a���}�z�;���M�1�yi�
Sf
8e�Vt���g7�0�´-�w��'r�+,����$׍+J֖�r�Ѣ��i�췪��܂�᭧E���Ư�s��/���Iv�H��j]0��쥣8�8䭱HÌ�7orn�vl�1�`�~�Gt,zeM�6�x�0%]\�>pb����O�819?�+N>b=.���:��%$m!A3��
��۫�pM��b�%�j��VK�Н'SY7��j��uwc:8J<.�s}�K��7����/j��C&�/q���s�P�{����	��@�'�sʣl::s&L'2b�wm�h4�$$:R���8N����G(���k:���
�9�'����u���ZDC)�Q�n^PBf@�t�l�KB2�ӆ�kOs^٭��jYD�YJ�!�[����aѫ3w/E!M�T��6d�t��ܚ���ӭ�v��t!��8jv�+A'-���7.L!a3h�˚[��=u��Ce�3Nfǁl+l+zBW.P��-�iQ����"�2<��/5,#7e]�9�d���'ܙ��k��L��Ƅ�1�X��L�uj����0�m�u��Y�����R�r�����2�M-C^a�m�x ��.�kk,sFRK6�ܼ�Y�.�cF��eb&�!�T�0m۝����o���3]�[ys3�ܬ-�w2�c��&]æ�]nJL&@f�2K�Z�B2�U�ys�@�Iޣ���͵�<�Q�QO��Ҹ]�{��A����)�7v�[���i��!i�d�7E��{C ����\4����f,��,9���3]г���b����"a�����;)��V�K�����f�i2�ѳel�D).RcK�[Wes,+ǩ�%�U���l�.�rWKՆc�"�t�B��,�7u�l�ŷ�<e)5U����n��b�։g�r�m�7�{F^�g��:�{��ᗮ�ݡ��v�Ҷ�hǕr^$��,�g{�Y��l��l,(ᇎ4aMY<t��Y�u�Oh��	(�4�(鄛$øj�4YT=.�i:U���eI��Y��H�e���WL�M�P�Q/fn�9r�Ӫ��$Y��O,���kHҞ*H���f�2�7BK���]1I�Ӹ��z#�3/�W	���2'ӵ��4Z�`��s���T:зv��,��J4-��=2���}���>��V��b���P.u�\��xx{�"gqm�9B��/���?:���4�z�$���p՗s�M���loir�xmU]��1A2Z�Rx��z��;*�u�T\*!o��Y��6��^>e�=&��/�c�
�����"�D]�6���T�[V�F��服���P%�J%�����+^����U����U�̐`X������qO`|b�++F�1O��\5rw]8pt'lP���������3��ck�b�W5�Bn�Y��a�,D2�d̓��HM7p�k@uo
��*P�
��h�rG�U�7á��Ok-PB�n���Q��๥���r-Ȋ�Ӳk�ʃ%�}�C�ۋ4f�,�뿱-��-qkZ���ԃ&��)+��l���Z�ُJy�����0ԉ^���aը�gQ�6N5��5
����D��"�v��YY�keFՇ\B9,֠�w���]!����?R�Տ#���-ٴ�l[�6��v�m�z̉�Re��ԛ��UTI�5F���r�>�g��g�8g�8ghμ�s�y���;!�:���B$#7h�l3V�[��F�U�FVfn=�np:�ĠΠ�v՚ܘ�jf���d�/5��8v��L1�$vl���y!*�.��U�,��m�	���	��e�*uhe�� �=[2.ͅf����ّ=W�̕��4ʻ�ۧ�<އ��*�E�Z��0�+4�Z��������;�	����w��	ܻ�J˗�g"�xr��Im�*7�+�o*�ڂ�&�Ư&ߣ�r�)�O&��b�7Y�#E��� ����lb.��3 4��t>��vN�;$�M�Q��1�TY����Bjm�Q��,�Z~+��y��1���ջJd0�G7,���̻���È�j����V�T�q[�"Zw�:�V«��.�*���pc������y��Hx�v.���1wf򲒼C)J�⑔�/	�H�	���o9�F�J�XiJG2�MX�� Cw�l�d���� ��
:Y[.M($[X.�w��Z�A:8S���mZU�hĮ��	�Z*TL<e|*k���3�.�v³��G�^�R�	�oI	�)&�c����0�rB�mL��a���^aX���+Ȧ�F�m�n����{�Zv3(6���n�"�K97���i�X�(���]��*8�s[��Crz��x$��_8,gN[�< ��>�IrF���W��aF����u���ƍ�]Y�3[e��ջ�E���Xz�|]�B�+c-��×C�`2���t��έh�)��!cW;L����������A��3�tT�g1�}Tu�09[�:ū�y���� Z關XC�bӌG��G����vYi���~T&m_'��]�������<��k�;b��<�PF�;�1z��� ↻����g@��Wm19b��*0���7V�9ݣ��i�,e�Q�',]�$
�0m��p'��!ڥ�+w*Ujar�6�AVV���<t���ۧ �8��t@�^�����9���\Soe�=�5ݢ����ˮ��X֍�����V9]�bs��P=⭞�!�������7C]�	��2�Ua;�C�ॷY��D�h0��9&@�LO�`�a�';f�̩��c��6������)�e ���lI�t��2J�n�+U��;xuf�"黗�ﾹ�k��N�>'tIl*����W������Jc`ӆ����M�!l@�Sc���5�e�$� rf���)ķ{�6��y0үN�ie�f�nϲJ�O����wl5����x�T���X-v�a�p�W��8%v�`�/�j�o[D�
�޲Ĵ�T9�ǘ�w�X���w;�B�h~̉�����ҝ����-�-��
J�2��l6.r��9Rma[i�àթ�u�r�f̛��=��9�Pw����+�V0kuYz�b��ʔ��x�=D��A[ڴt]�f��F`�iݍ��X��!���LژT�0��,n�UvtLSS2b�����&�n��5�-�ʊ(��3l^���������ɝyՀ�����s����Kb�V'݃����e�Ib<b{b�jn�Xt&qʶ$U��9��7:�Wh�LX��SJ�Al2e>�Q�r^!35�k�0�l�}��;/F����@{��C���q엥e�R��I(�5w��c�g��l�HJY{|��u�ګ��먵"Ɔ4�ۛcM�S�T0&t��s	�)��CY\6]��C[�]���껀��s2��U��M��n�2Q��Qu$�4UQz��1E��Vp+0�.�nx��x��9�\t�vv3�Ք�KTз2� �J̤^;|R��C�r��V��x^!��ەuc7sNc�V�s9�j�'sLYW[�smHYA�����Ki�c��*`R�HK�F�*�Ä��9��D��&R��F��^��ֺ�r�Y���E��	��U��NQ�M����&Ǘ�*ɝ&
j�t�b��"��r\6�d]L[0�F�Q,5�Gv5�T0*�ݴ����C��hx^!��hym���y��Q�HȲyίu��K2������|���l�R��Bl7��,��w���7���.\b�>q��ˌ{�|q��S�>8Ĉc�87�ً���c0��N0�q����hMCâUR���v��Ԩ�W��`ۺ{�)�61��&p�Zx�Q+����$*K�굓��fNL:*�U�I׋F�c1��T�%�*������*^êY71��C&μ��� ��bU�й����̂��cka�R�11˦�B���3l&!�8��d�B
�vx�\.�����5,���P�+Se�7����l�颚N�'h��)��	�	4!�)��t��@N	�uj��l��Y�G5��px�o1PNUJK��N�-�J����.�9��0r�rMTM�����I�Y{h+]�6[����twz^l�j�($]�ܺ4"4�R��j�ff����[FlV!ۗ��'�i�r���_pq�"Q�*c����	�2�;�A�����aR��Z�QuV�6ȩ���Ū4*��uoeKw����cf�"j���9x�bt��4��6����I�����*jw9�������
�����]��+.]�sf�02�+�F�L�Tn�8���6b�q���j��n�/q�6l�tk��$(��NU��w"�Xv��Ѵ�u]M7�=���YB�5�*���tCf�<#ޓPd�5�n�w2��f�������M�����ӇOl�"[�]��T����$���S�̷4m=���P|Ѽבl�U5p��_���1P�È�pb��T�0>��T]��9p�h���z�NIY�2[�a(<�!��TvTic��U*%
X�V7�+o4I���b�,����C7i,�T�;�1qm��{WE�5n�`�2�Xq]�t���L�̛R�[D[�SBy�h��̜2�m�'����g+���Φ�W���6B�Z�w�:�Ɔ	}��)���;}�o���NV�Bpɘ�{��[T�ON�3M5]]��BO��r�zpH�XK)S����*��薬]8 ���1�:]�BuĖMK�c���gm�Fݽ�z�t/gi�h�E:��=�����a�G�`�Xp�@)��o+CN�z��iOo�_�;�;8W�T��Vt �(N1�8��`�֓������T�ťd!��v0VܚA�&�e�Ro�[b0SU��u(H�
k�W����(�Q]<`�ӵ���|_	\NU�+S�<xr�^ޡN���B���ʍ�ztP�wq��=�+B�\s�ێŴ0Z�^�@tDf]��r̕K@�-�Iz�8;�ڶ�lQ�	hwbs;�Λu���Cvej�bh���ˑ�r[
�f)n���^�����oպ�y��\hяM����r�j)[�
�x�_PZ����,es�Cv�(���ɡ1�5d��#�R4���QQ���ߐ��s�,�]ϑ��ʌ�`�X3V��Vt-�銳lk]mhةm���y���V[����T蛴iPD}sS+�g�����轨_!�,�:+U�'����EN��NXf	�ٍ�;\o��AZ{�Ch[��7��+��p���'N\�C�N�!K�n)�J��r�2��E�շ�-UV�8
k�|�;,�G�ݛ�����iKF�����d�v�K�[��UnR�U��/)L:�t�80Yڇ��CwO�J0���u�=*��d���D}�t���$�D�2O��ӧ�I$��Y�G��z:h�eQ��Y�,�3Gĳ���E�>��iq�E�h�����A��Z	�����&1���v��nr�n�Y��%���,��$��e�Y{{m������I$�I$�Ym�ݻym���I}}v���d�I$�I$��$�$�I$�I$�I$���,���\�I$�I$�I$�I$�I$�I$�I$�Y}}}l�I$�I$�I$�I$�K,��,�H  ��t     ����,��I/���,�I}e��m�I/$��I%���,��I$��I$��I$�/�I$��^I$��$�$�RYv��/l��,�I{e�Yd�Kl��,�Im�Yr�$��e�Y$��,�s�m��K�m��I$�%�Ym��m�Ye��m���/$�I~�\�I)$�I%$�K��]��,�I%۷.^���$�I$�I$�Kl��,�I$�I$�nݶ�$�I$�I$�I$�I)$�I$�I$�I$�[m��$�I$�I$�I$��Ye�I$�I$�n߯��l�I$�I$�I$�I$�I$�I$�I$���$���I$�I$�I$���m�������e�I$��,��$��e�Y$��,��$�[e�YrI%�]�r�d?����I,��,�I%�Ye�I.����������ٙ��30ff��O�����Iv�,��$�l��,�Iv����h�V�f�33�ffl�����}�l��ٙ�ٙ�>�m� ~� � �O�G�?NO����n`;ff`;ff`6���m�����ml�I�ܻ��ٙ����}�ff`6���m�����m��I,�ww��m��I$��%�$���}�ޞG�?P��O�ff`>�30ffa��m��Ye�K�m��9�  ���������}�9? y �� /oٙ����x^�w�ffl��ٙ��3-��-�������]��-����{���33      {������  yn��      n�t   ������      9y�    ��  f��        �3>���         ��� �33 6����m�K��Ŗ�m��Ye�Y$��,��-�۽�{� o��m�I$�I$�I$�I$�Iv��m�I$�I$�I$�I$������m�����I?�r��߭�m��I$�I.I$��I$��K�n�l��,��=�m���$�䷬P�������_	u]���6�It�/($�$�F�>0�7y8t�UUB6����e��[ff`?�H���9�v�������xgu�{w������p���z8�b�9s�ҫr�X��1�]p��xVΜ�k�ݫ��+>��>���C��c��+y6-�<��{+R&
e�#�ؽ��X��!<�&�Ի���_N]�W&�[ĥ<P�V���D^=q���f��MNُj�?*�>�Y/I��jl�y�0{0%�a�X��'�XJS�x���]a���h�:�V�n�C
��M���i�Y���JKu%�FkK��c��w�rO�*�!�T�Runguv\V�v�o��B���W�e*OS��5�7��`����T4G{۶:x��u<��ڽ(CudS͆��6��m��7
,P��;��ki��t���>�H���Û5o7H�$&H�[�uUo �U�R�3x�8lm�m���{���^�p�NV�T
�{Ó�h���Ⱦ�[T��o�������1��ɚ��F�^h�Վ��t*g�RK�<6�7./�Ů,�uŤV(p�=�:�8��r�qa�nսFu���k�⹬�a�7/cC3�l������gXب7�VQd�N�P-���3wX���-�1P�X�h�F0e[�������'��҄��;���bnoJ�	XwfS�Z�s��kR�5X���g\Ж�6�Xꊰ�L���;M�[KW2Ҥ�[�Yy+j��m���p�W�nm�G��V��rvۛU�|P���G����ʃV�(hK�*�	;SER�̔m�*[ pr�����q�v9�&������`�ܞ��3��k��͈�r3س�Κ��Zu��v���8u����1�8��89�K���
��Ud��o�htr���z����a�Q�&"�UKn&4�Sn�.Uh�8�#�¶����.ToQ�m�ӡ+��j�0�TDinҫ�����k���dR��^����8�N���΢�V�����;r֊�Ϩ��(���nvцKv1�Y�H�*[�{�e�A�.��Z�z��\�KgB&�&��t����mލ���m���H�T�5�b��:�띻W$�z)��s�<{%D� ��]��V�p^��=ձ�iI�1��Y4�;-�V]M������=*��0�䶥�Y��QmX��2Y����_>�E:���ov�[��y�+*�K�5Iogvf��MV�YQ���%�(��3�o
��4�HZ��1j��Xi�K�$��( ��B�9ʦ�8�U+��n�]�;Z�q��v���(�2�F$5U� (*�{��澡�Ko��o�V:�2}�m�����AN��ࠛΫ6��`V���(gm���In*؞nw���E,풻36��t��zZ���6u�g�15�{�i绳�͚��]�}�)Y�����>ךÝ�^�Kc���Yۓ�_�k�����U���Gg�^K��C�Z`]�:��x{S�@�������h&V��9�a��`��wfeV��w4`��dlȝ����6���[*���"����m�,�s�q�֤Y�2��	Uqd�;/L��b��:��h�^QV��{��w2�K3Bࣉ�ϭ���wjo�k�I��+qu��}�e�W ��^�P�ĩr����ߎɓu˕�V�t���R��܍�y��j/Z֩r$��5R��+�b�a"�-)b��Κ ]ۻ��d���f����R��J�G+���`����l����X���6.wY�����Jz ����^�����U݅E߹�uc9��A:�7\���Uݔ�;ؑ��&����U6E���q*+5eGv �؎���mUm&���Ѽ����CrR�]V�1��J��%j37i��伖�g�Zl�)V�o�f0�%�1&��X�e�tYN�j�I�c��뱢�J�i�|�pWZ�'����ï﷖I�M��U*��}�=s/9��voj\�.M1g<�A(�Ǘ����W������U
P­��	T�ʾ����W�v
gu=!775a�S��M��i��͇F�v/�.�@�S��^oj&Λ�>�*^>�r�9��e<I=�BQ��n+d&$���W�x���'�s����ki�����]�ĵ���ڴ��V�	��뻸��Y�a,�RE���iS�K�8j���WwmA����<�M򱏲vG����A`ί*���;5��1UцE��<:�Y��Z����-8n�w���GC��.O�߮)PWPo	���l�1����l7T��˓k�)VI;7T���r�k}�;h�n���q�.w���γ[=X�N�nUK"ى��Y�%e
�4s�<2��t�}��˾��_�٪9Wz�SN�N������y0pyn���Z�-n�ڮ���ͯ70z�7X^"<]21�q�?<�{5r=��I���d�TU*����f$���Po4�U���A�����r\2�,l�ؘ���K9^R�Q��n�Y��S�MJ�	N�hNF���ŉj�\���)6��Ң��4;ݳO��[����7��^A��P'^g�dh��I|��a�J���%��7&�����]�)���-�`5-��k!��^������0�C�/`޷�a�v�+�˹Y���]2�ܷ�e�sw$��{@݌K��_K���7�Q���Ԫ�H�a���b^[7��)t��	ŕ�u-�w�s��wۆ�x�fi�)�p鹔�(����Q��;{ۤU(���e�;n�A݈q��e�ﱄ���4��14�s"Ys�P��k�2)�f��Kn�=y/�N{��u��Vu��|��ԕ�ڦ�*��� �ѧj�-V�E��r�N��z�XA�<���e�Gb[�F��:���!�^K�"�����,��^�W#ھm�:���d�\������>W��n�Ƅ�WU�XM�4ƛh�oNղ��S��hT��س�ټr�*�eB�L�͚�U�C�1/7��˛T�U]�M�1�@�6�-�X�Se��_*��׼OK�2vv4)���Y�X�L�0^E8XժՍ»]�@�٥R��D�R�ީ@����a���Hb�b�1w��	+����g�L���ٴ;���V�D�}�%;[b�l�<ٗ.�:hA�r�X,�I��4���o�͛�4�$u�dh��g{�9�5RR.U-�F5�aZ���Fn��7��1sS�c4՝K��1C���D;�S��|�[��,˪Uu:r�bT�umP�NȌw��ji�zz����r�k��叱�غ����
��ڪ�t��فQ�����ż��H�=��({2��Q�����1b�,�QvH<�|��E�����}��[[��,�,U�J�"+W��z%u��#-��A[lk��;PiM�ӆ�af���l�·neR����b���W=#��u}�6�D��-�:��	`���%�T:��{�J�3u;�Mv���+��u"i8��r3V'�"�Z�
���k�'��șe���1�{"��.���~��M�uٲ���^Ќ��ۚ:��3bjv�Y��\�:vf�������%Yݾe|�y��Z�ޤ�f�u*Kݻ�*��F��O8&WR��z�썴��y�IjbJ�B	�%B���4KHT�[*�f�����Q㦜F��k4��d��ju��-�{�r��^��
u���fN����Y����1�l����0]U��-�T���{˸�u�u��6!��*�ٝ5#;:q;��U9.���ɳYL2�i�&*�%%!{�b�A�mثd�].�P�|�䋹��g�oxZp�W�Xf�]w�]��b�35�����إQ�cn��ܵie��t"��F��~��[��&�Z�(D�<rlm$�`�6�R�مf<�O��m���Z��}V�Nj	S��Ӑәü�I\���M"\��j�kW�f���������98ڑp�mm�6R{.���n�U;�:�su�)Ua]B�D�=R�F�nP�yΗv�N;�=��-k��[''g$�r��{.Э�o�*C��=u�N'�#s�Sn&ʬ�@�+�jP)�siXV�Z��_}O���̦Ƞ������kuN��m�i麊	 ZcJ�o<�UFd�Fc��X�u�3�팳/�;:S��8n&6 ���1��q���uf0��U��9�2��U��;n��=j�{��m4���R����k�gf.�D�xET2aTS"�A�S�)�c㘌�.�ͬ�s��v�6�iQ]�l��a1�<�,�)Ø�
���p=��i�n1�u��)5��s-ދUk�K2"�J���bm�����x*X4�G�3��5�k]�N˒K��s�J���!'Q@�+�
CH�[���w�֋q�b�T�C����� ��9�Uŧ�Xc$�-�/nf5�r��*�*���W�ฐ�{Vw�����}%\ؠB|�J^1ypZz6��*�펾����jQ+�F���p��W�aWx:�h��F5rVMP�|�S��s�+�Kn�:���󟭒�����,j��)�0�K]K{�կ#,��{֬%{�o��]z�u��ы7{Q��i�ދ**��Pռ3��:.S�N�|j�}�r]c��{(Ȓ��T;F�If����zk��6α��@��Wz�}X��0�Wy}��kE'�z���8qO<�`�}�l"��d�R,��4�\�����V�s�X���tUkyT�r�]���%E�U)���"�qf�ESɛ��ξ[����7�m_qAg7�1�Z���VÆp��y%u���f��
��-�S��E���\�Ů�N28Սe��Pl˄Ʊ7�=�Ie��|��jr�K�*6��U���9|���z�_��/Ouc9a:������m
t�	W��c����:%�ޮ���r�G.\�En��f��*:��\�k�ȼ{��|�vj�DG����a�J�1��ИWg���ʅ�u�D]6�ᴡ{\�5���������ܹa���#V#�elȺ�i��ݣ�x�xd�rC��du�˝ח<����OwJ��iN��뉃,7��)l�>��ө68�ҿ-��r�DxVeR��bjr��C:_bzxm�[�#���
}��l$DR�飝���w��IR��Q��d����ۚ5���F�u^�ah�v;�x���RYTY���c��\���-�!Sл/��L!��ԺG�C�<C�q���}�Y6��}�O@Y+ٺ��sR�Ul��jхPd�
�r����}�G7���!�ͬ�i�Y¡��K���ȕ~bHDH�@᳂^i=$��0c����v!��ү�D���M����}��ֺ�99�oe�N,="�<w�.=��mn=�����N�<��X�+��]����1!u)Tga:GN Q�+5���yk�+�����v����FN��)d���B��k
zNs}[��GT�g+ ��q��[�j�cE�p?�>�'6x>��B�>��_`{�'Kh�8����fV�}��vjz��$�t��yl�Y�¨ZZE���u�N�*�t�tJP��l�T���u���lf��J�9�2X����!/�v^bo��*�oMT�p-�����Ѳ��;I.�C�&��2�Y5rI��5&�P����
�"5��]�[
�T�ݰ�V���d��K�bm�rgU��;�vm%�U!��(Ԝģj�L�2��G.Eh�ɔ]d�iF��wiٝ�R��^���~w���?���0?�̓`}Ct�6e��W2��y��
������
��1�g�Y��Z]tv���o3��ť��[��57Bn����*2,s%��x���a;&�`�W��u��|�\Ǳ�7��[�,a�A�ѩ#��01�suqi��N٣��Gr�h�� 8h�2�gb$;h������8��7ֹ���p[���%9���R�y6`��b���Π\�
,$�	k9pZ嫪eI�u���oAvt,;Ԣ6,�.��'vMO����e`�1[e�~�n�ۈ�a=z	l��o�j#Ft.;��F�4��MM�c��sO-l�l;j�DN�����7�æ�@k��4u�d��[��՛֮�uv��['$��@�w|�-e��|�?�e�ϳn[�qs�q*Xkz�Y��u����jU��n^hv*LA�Ps_ܲ�w��ں+��fp��sb��Hk��:���oI���u1U��%��f�d|]s�#74e�nM��M捤�UQP͢(��*�Tӕ�)��u"�7ZRY_No�w�]w�a/�F1�����q���q�b�.K���9+ѫpވɗŴqp��ƚ�F6j�Y����sQ�pJ� ��J��'�;P�E-oM�r���n��]ݵ��n܆�$X�U�.H!x��R�R��H�Y.o9v7�l���6�����Hh��(��nV�����X6�0��g>�C+��%�F����|�\+�5+��k�hT��=uӠ�N����8q�N�+�zӥr�b�u�w2�]j���K�*����^���;�-�髞ؚoN�]P�]�c��<�i�$"�|91�i��x�발7��oF{�s�+�uT�s�_X�Ջ�4�X���J,��^�/b�����j�jN�Ι���];�[�o2w�p�L�3�Pk3��2��P�SE�>�ܭ"o�q�X����d�2����w�݌uN��e	��$�RLc-������k᭖�t7�.��C��
RͮWj$�RU/3����ql�Ӫ��U��#K_u��U5�u6ON��:����ۼz���4M�r��g��f&���vj�P92ʗb�)����8��	�ә1���Sb�]Ns���8���81�=��%/�)u�c{;��T�qU}R1y$��$�j<DZ��
��UJ��쇃Ǒ��x��T�+x��v�ͫ�mmud,���wE0��J����4�X�b�V7A_��Su��셺S��v�D%f���U�AYl�J��a��qg�7ez��8|QB��q�Ji��[x$9���+��SR��ڰÜ�u�-Fj�nj�㋁��F�o[U�iؖ9mu�Z��7�2�uV�(���f*W�u�����4olZ��\7�RF+������Q9p�X�g]�Y��]��yu7��������|,q��z1��jB���|��/s�rV�p����gCC=�u_����iҼ]b�܎��[qpy[���m��,��v֒3$�,��������[��]*[�#𓧞�������C3��8��k)Q1�w!��g�]����K���'�5�"�1�]{(�����wSPe,/-�|w�P��7�G���v�Ano�_v��}��HF�!�6��eM'Mlm�{8'l]��;�p�;��r�s���	�e�t��##ف�Vn]�O)-Y�)�%���:����	�|\�j�AZ�▹��U'��Ɇ*�Ô��{N���+��E��`���f��r�s�n��y������nr]@����!��ʻ2���fq�v��[t��L�ve�z"ޔl��9oˎ
h>�m�*��q�J��L�UI �9�Z�-P�I�����G���Wh��4k���'	���q*9�mvt��;�,�u��ӭZ��U�eC�����>�=���v��"����o2�K�:� �nȫ�75Xu[��;b���b�2��.�Y/���9�.�c���{����� �!��Y��&{3�*"%
������^)�a�r�g��uV�R��:�C�h�{���ȶC���j��V⼀��.\��oS��GO�d�q��&]�zp��趫K
Ȃڮ׽j��p��n�ܓr����l����+y��f˯T{�$��;2�p^�&�t�%�ܴ2j�y�Dc�ډ&N���8��++|p�m#=��N*2���<�pUYH�5���b~Ⱥa&z��ԞQ��j+XWYp,<�j����p�i5������m��A��k
�ǳC���N���S����6�_R�������s4����Ə'��/y��T��R�w�Z����!Ӑ�|�.a+sgVp3�]�84ڡ���<��'fW}"��r���r�� ���SG����o1j+��JR����!�]gN�Ή��б��v���ɹ�N�D���Æ��*I�;6j�19sL��N��t��
��^�=�s�F��������d�
��
�=�ՠ޺�E���k5Yk �ʔ�R_
��)����9q�չZ�R���È�͸�s�/'�)���t�8-T��$�>����S�V �ڤ��:f�Y���F�+5�0��� �U�2�h8���NU�A5���6�!����ʓR�޶Q��_J�n�8���/2��V��K��J�W�x�]�vr,:�I�2ڧ.�|�ud��� �sh���S�av�OM�j{���m��"��z7ެ)W
���-:9�PjV�ƣ؝�L���
��9O썂C���z����u��!���	Q#��i�0�Av�Mꝴ�$M���R]AYT�q���_WnMn�mn���k���OvH���X���D؃����%�c��$xѼ�0g�ۨ�;�����m���9�YaP�b��_RΜwx���\�N2)]��c95���'-&J#*_Wo4r��=Oa����|�]��"0q�;�2FѤn7׽��٢�s�3���)ґ�q^��NL�cv��C,;�j(��a	�[q��o�Y�Z{��s�F�9a�|��o�.�&6��[s/�P�nF:��a�N�E����&��Š��Ӿ��b��T�ټ�[�d-1�K�#pZg�⏓12���eM0�6�zL;��a�A^�G+�s��{U�8�+���7��2d{/f�e݌s�A�;m^ɖ���[.��n�ы̇�_8�l{K��S�z���EZ6˩��՜��j���OMw~�}�C8[8���;�v��j�K�]����S���sJ������]h�^�˷�L��t8M�^�}d.ߺZT�I�"�Y�ᡱ	���ǵ�UÙSu@��s}N�S�M�7.�'��+tC�9P��L39��bw'E�Z]
1�h�����(��JӼ�����Y�9Y���kB:׺���|�ov���Un��C�#��Ԗ+�X�Nt���YBA�:ox*]�֊P��O!����.�+�Zx�:�L\6�M�x���rI:T�/����آ��fr��n� ��T�F�9�Z	7;2qG���Z PWg;4�5�p��4��3����k=o����N�n�?i�v��Ūv.'��+�
e]���J߸��T[�كV<�ͽ��ә.^�N�S.�.�:H��,b�^���7�j[����*�R���']������ЮkxԪ�f�*hf�L��dv���\�4�7��.U0s�\1"-L�%�m�5(CW�Mw9�Ĝ��Ȍ!|a��R��L)Q
[Ulr���6k[�y�j��R�7�h�ձ{e��`���4�J�d��a�X(�3GWlt�3--1ޱu�=3I�#7oN��z�Z� ����t�)rGk��Cm_�[e��Ý-u���%+L�Ѫ��sp��5܀�����,o�7^V4Z�>�uIjls���ʣ�9���Z9�j4q�	0�V�-�� +��tG+P�k���ǷۨT##�b`��[T�9]���ڬN�����"c��;�O���f�v��Cx:9E�:�qgn���Z�h06޹OL��S*�^�q{�1�V��!�zֲ��S�#�F�0]f�*�YLj�.��y�h��n�����le�Aj�ڕ�h��j���y|fj��+9��MW"�.��%?1�k�|�^*(0��֛�U;{$T6���;V�3���^�1�.�.���;V�{Z�0\��;L��Tł�¦l�Z�;���c�����\ә�g�ug��
��J��j���.�-[K0.���/0�j��1�z���+N�uzʁ���	����Ko�m�7qK�[#g��>��]ŲL���Hl�A'�M�S���c�nߥ�Z.�&��'��*d�|E�u��5|3MtȮ���{�ΐ�)��"9��7�_v,��֢�k��f5��:�-=��������'�i�g[ݮ���u��[�S�������Y}�[O�X-6]+}՝�9���}�eF�'��'z�a|����>�oAK�Yq\�X���8��]�T/�v�r��͛��0�Z�OW�x2����;�Fj�Ж���z8o����[΃E��樯]Q����0)g��^�Co�y���'�$�o�{gz�;[��?�	�%1r�;�\Wi3��=��.�\s�(TR�v�,J��ǩ�EZ�,�Xzʸ��*kB�
V��i���8�V����wta�{�{�����}���SI*#i^v�ʙ��W)w[Ѕ�:���X$(#3u@�|�\�.5�jq���N$�&�6-
�Y�
}xHc';�c�ؼG�2��Q{A���@���$CX����/1�*����@���E/2���kwb\peԨy�7������gx_E�n��������o;��U��
dM��]J�`��'T/.7V#ӤSB"�cl4�����LR�M�,��_�|��[8']�NL��Xgq��`��pmJ���d8	�k_^��ۇ-rz���kY�ʊ}M�y�^��f^�y�V�ĻVA�6P��7^tw�S�5��|�Sd�D8���N�5:��;�ì���0uP{Z!Vv�y�hL�����ꕝ���k$C-ξ�V�'�VG�m��Ȧګ!`=4�t��+N����pH�#�<#����=HgZ"J���BtV���Њ�-D�4��}}-���t�[���4\;U/���B�����7�;�Es+L��Q�aQϩ%o��OmI��n��"MŹ}��g�S���R�}yr�5���$���=|���}y́��飡o[ZC͖�`�v�G��d�	\6)�!�*�eI���%l�]\_0&-�R�k��p��(��n���V�ϱoX/0�ci�t�3wi΃�B8j?�hnК��
m��Zhh��,պ���7x�R�5%CY���+ea��j)9�ᘕ�]0V��^j�C��*��z�n�+[��Qce��{t�+/%�=��ے��`�u
b_>�N�:��o������:�s8ҡSzӼw�0�
ծK��]����M8�ֳ����2�u<zcԢ�/����f�vK�'L��%6�e��y��Nb�6��}����&���><����̫5��'��^8t��Wݩǟ_]�d3B�Z�=l;ɵ���l�o�����7�R���K��լ^'U���a�2�h�؝�oziGb��&�_���xx ���6���f�V͍��OK���?�l�r�o�I9�s��䤒I%�~�������d�����m˗.I$�[-��l�v��d�K�<�N\��go}�6��m�I~��}�ۀ]��=�wA��N09� �������������������g�� Lu;cw�؈��a(�Ʒ���n^�]�$2y��&3Kc�EuZ�ʦ�ߏ��\��#k.���
;#�Ŝ;������<�g�T���V$�#/�k�U�nouV`��*��Z�*�2�iBIa�ꕣ0q)x�ќ^uU�P�=399z[���҅DN*��܄&+�T�<zpJ�o��拑do���ʍe'A��lz�Lg��}��;Z:`��x�w\;�Ӊ��if��K�J�r�v��*u�ǜ���˳��.�]�J}*J;TFU}����9.Y��L�)�����*��o�Gz��I���{s�+���ro����dm�y��uW�w�M+qb27뻶�S�i���\ıS���}{K-M�w�ͭ�י-'(�xN�&�W�ۙ�T�+�Q�7��W�ֽ� ������ڵ�sdy9ח%�����E�緳�m�&���Lн�`�UU~H�N��+`bS�^�b�ٓ9G�`R��E��'wu�3.�5&Nְ]�7�8��`���gL�V:�4��pWc
�ګ��J�)��[cgGչJX�rNӧ�U�a٤��)(��o��ͷb���^��	�DO������6s�����k:�M�+��@Y��a���$�o]�.�5w�1Tb�VG���d��5�\�מ��Zv��dT�Pl�%�L�����v�fј���,7�#�HȸoEN�*�%PtgaWzŋ	AJBYWʆU�j%y3hغa'��*��n��U��ݧC)�ċ(�8�()ܱwv.�H��y;�(ٝ�1+���n�h3a��f�K�*�,q*��p����.����ؑ��d�b��4ʕ�DT�	,�	�Q��C#���S��/¶�Тr��P�
ahK� &�rlux#Ң��Aw�W��%�wK�~X��9-�yM2Px�\�M˶F:rX�w��餓����lSiV�j�زgsf�$���P�Zt�W��h� ��F('1T�+"�Z�$�h��A^gR8x��<�� �;�|��[Xg�ly($��2�a�:*��R�8FG 	[Ǔ�e���`LJ13ɋ���T6�,�֦ZB�Mh�i=��x��̆࣡[��`ؗ)! �̅��Ӆ�U�'����A�y�k�UG��|޶��!��0(\*�\U�Y1ژ�vX�;uF��Z���7��C��K�n_�+@�(�I32�,����hU�ř���!���`��!��`���(`c� ��0hJ0��4[�{9�n��1�Ik����
��J�5[w��wʉ
]G�F]��)l�h�DkZ|���28��:�v��u>�Y�ܳ�ռ�Q�qY���71�ǿO��Ӟgӯ��� �H��:����/��c��ջ0�/�]�0��1���� <k0�ۑ|�h���1���X��D0��C0��%9�f�+غ��R�4�,�P8�A�Fl,�_�S��̼��Y(ܑ�/��Ih�ew_y�\ւ��c�< b� ���B��$��a���2,K�>4EZr�>��}G�Ðhjǳ���E
�Y��Ra����Úd�z;�}SqPz "


&G4���c�h�r��|p�Dѱ +8P��)oՕ̢G���ͳ�p�8s���:]=����0��*>Ԋ���C'F�f$�)C��8�]݊���6ԫ�H��x��ݣkcL���417ut/��u4cy�ht�P�Ni���1s�3M�fI��~{�}c|�ջ�rm��)��&rok9l��nM�ML�|�rc�	+m��﫿\��;�R�d�S�@�<92g�R)�P�cwj+猪 �c(P�E�� �4LC�k3I���/|�I�n�~I�C^�M% p�I�A�������'>�Є@��$�P��{�S�H���m,I��@�H`�"���yE�_F�b^�0�O�H�1!4P@8P��������h��7P͏�(B
�)�F����q��n��������)�즲KA}�k�k��0\!���
��!DB=��lA�{Bᔤ��ZP��l�Ip�H栢��k���	��fj�4V��ڮA�"{�����i�w�Q(p�uDm:o]�������91@��3bAI�>IvN��n�r�M�<�:����m�V��t��'0���x*��OI��0�e�sd�v�M\q=V�h��> ��	��nMŜ�mG��K��P:t� ��	��:f��G�ɸ�QH�,�&&q��M'	�������
_f�@�A29� �h5��*0�l�z�=�!ǧ$E��R@e|Ih�5ԟC��U���0�$�`��l"�H@���6h߶�6Ǫ{r�h�I$r���8H]��ums�%�L��ҚJ@�~ �ǈ3��^ץ�$��s�9H!Ɖ#Ĕ`��r���Fb��%y�L�� �nl�ad)��ǉ-�Ȓ�����o�D�������ɊF��UcnTG��[��P�L(| �NR �	@��ǘ����d�`��pwC���x��֌��/���H�{γ9e
Yz�����V��[T{z�T[��,�4@�{wy��'z߄A�'�6M�L�Q�5��"�)�l�4TL���_K4`p���*����j^�`F����V]\պ�u���}��9�xRVC"K��!�f�@���2鬒�DI�Ŏ#Y�#[�O�s_rb�(�$'>E"P�@��aG�U�>�>��쨮N��b�1���0���M��[�#�b����G&����+�6���p��n��q�,�ds4��9h�b�<	!��	�H0(� EY� e���(��O9$����b�`$��|��H@��O�4F�9Y��ڙJ� M�ŎA�b�>�M��!�!A� �s��s@j�}A� BEx�0NQE@���_E��<Ky���$Y%�NQ�["�u�!o�^�2���q�Ҡm��6�o�����'���\� ���W�E�ڊ�:T�����/~ꮜ��4넄(^`�0P���!!
# B^����U"��t���p:m�z�彭L�7�4d�Z�W>P�j�ީ��(�U7��p���X'�6�}A"�	0,{$��A�@X�a������KE"��g��|ȹ�fl��9f�)�>r����$��̀}�w1����> h�����
B�dbD��5��/b�N��+��{m�KA}'Ɩ8�0r�!9��C�%՟z}�T���j�	x��V�����I�{m^���z� ω�Dy�0�ǉ)6�Y���[�Q�|X�$��i@I�P���>�EC҈Z��m,����	����Lr������Y�{��6���FB�� �KD�y� E9�7�U%���*"��5�l�E!�B�Ğ(��I$ߥ�t�/~E"P{u^�y�	���5̉�Au������E���s6x�^M�����3p���	p�A	SݒF�^��R�I/N��4^�Ng��B��v=���UG�V���lrTn�{7\���E�Wj�F�h�k2�A��Z�"\�%r��{
!�5P剈r����b!��)����%s�5n�� p�4h��NQE@��D#Y���/��o��K��đ��94��4���s�:>E4�t3 �O�&S���Ih�A$�0���t��sb���2S�K����xr��@&Mm�ɿ��7�5\��Q<$0���8Pz�f0��}_LEL�1�b�d��G�T�'<�F�4�ϼ�'|�|%d�Q�*ӔQ��).���}���URf��A����$L/�x��8�d5�0�G�%f��e�	-�R�'�9!�oL�z�{M�k�W���DS��R+�X�+K^�S��Wqv�;F�4��n7��9h���t�6�}��@�vTu/S]	���nT�A��w���tk5/-�0�n��[v�Uvs��Us	y����m{X%$8��H&�e��k�O`�D3��������$0��KXi'���Ow���@| � �MD���8�0rd>���ż����oǒ��3�Sd�Q�,M$�9��1��}��1�Tl!"DxD!�~������KX�Q��v<4X�'(��D!��	#	5��ϗ^�ݫ��Rr���-��x��g��^��"�ts�Rpw��KE"#�A�)�3<}[r��&KL|��a&�P�L(�A�Fi�J.wۆ4#Qdy"D��)�=Md��fg=�yy�Q�P�z�b� ���hh!�};ki��w�A6�g)�8��N�%7��G�Z�]=W����p�!n�S�$6�v}�}R<OYs�0��
P#�UU�}����� ��XĶ.��z�XU�n���Q	����{��5����������7�3WklC�2-aR��UN�J(�O���Z '�Qb*ӔW�H����$G�k�F�м����^(s��,��8���ѣ��'\��8���A�H��P:'�i���4�<�����D��JH�h�l׽��N�^~�y�"G(r�U�"Ȳ;��N�\�%��`��g��4�#�|&�9�4�6�,YL��X�oV��Rk�	<h͇��T:�
�hP@�D!�4H�0! �h�ܽ)�ɨ�������'�,re8>��mO�N�^Ah���>(p�NI�&(u�~�qLG�Q�"o��a�����t��Uȭ"���r)�t�]�]#q����,�r�A�]��kM#��R����њ4p�� �Ɔ�Ѣ�V_�1<�����y�h[Նի�l*���SN��؊�u^�;]���)nj툷א5��^�p��-�D(�,�$0,ꈨ��~$��B�P;��✤hޫ�<�/+�F�)����KA��l�����UM|"E�HNX�D�� J�>(�0��'6_���0��E%�D��AE�h�#���x��χaN�I��K�1Vd
�}Sg#�|�u���)�$,�	���1�f0����ձ�,�I	�"0DҒ(�I-�4���j!�vLC�9�!�h�E!�B�4�Y^��}���wr�X�I��>B�>�H�y�}w��*Q�����M% v�$��`�ԯ�>�������b���C���֋��xҋX ����(�+%�nb�?4�����c
0p�*�Jc�����붛��;E���+�Z]�q͗��]�cY�ϝ���;k5�.�0#�D�e���7E�	�mj�ղI�P��ڊ��a�IY�V,�R��P(������`�0AC�� �A��M��}OPBu�P�Q% U!(a�8$q����Hz�$1��D}��a;��������Pj&_x�)G��qy��[Qq��Md��#�>4��h�D+����W&�f�'>H�6%g�(������}���{�2_�X�� �$F�(���<I�5Z_^���E���x�Uz������}������#e�L��x�-�au;;��ws[䐼H��JH���KA1�"�sriU%���E�V���6P�ݙ����)�"��mE��N����cU4�Y�CDxwq�	����j��Bś����R�B�՚��4�Q-�WJ�F5�(bVsU_�ѹb�!��ט�w�%u��%�2�Y�:j�������ҜXO�E~t8�9����?�k��'KQS�ZR�>K��x:�yWv�y��]mMD����#F�k��c��u;T��]��Wz;�9,�$����{��ݩo�y���0����f>"U�nǒ��M�c���*�I�N�А�[�G�+���/L�3o��~�թwd�EKlUB�r��H�Ӻ�͉���K�ыzI��KEEU{j^���9U�efEV;�6zvoWh1dz�=���X��)F�s���N�U��e�\���Ε�G�������LXƖ��*�딪��\��fu���[R�eeS�$x{z��{P$ӻ�䶷U,�۽�Ө��Oq�t�Fܬ6�>�e��T��箷1k��4-�[�UV�D}*�Œ��)<�I�d)M�)�C���R�$����]��k����fӴ4��b��#%O=ܡ� �s���������C|C�F�����|����G
���cY���%��c�i���#��;y��hA�81�
(PIK�n��l�I-��nݶ�����I$�RI%�~�^^^I$�I)$�H0`ѡ�� �ltA�vf`���3wt＿^�_�������� ���wt�����t��}��%���I{m۞[m�I%䗒CEt�'d�7���<`좝vB��eK��!�CV���uTK��Xr�8v�Ώv�j���P�����\{tsiΩ����ܚ���\��I�#�����Kx�mK�סꛋN����e�jڪ%P�e��7�3�Qn�[S���Ro�.u���nW�\��.[��۴�s�wW;(�k��aP[�6���yJ�����wēam'1���ҡd��5Y�t�R�^��kM:��`#u�WISk�	P���ϒ�rjӹ���D���:��xE�Yo��->�<[SN�[n���G�xgAǘ����cd��_S\�̊���z�`@�IxF��sk/D�]�������3��W:��(������Y�w+|�,���k_b�P�DU���ζ��~Ǝ�j��N>��*�CT�F�3�gf��@ͽ��h9�"�5�[Ó��'C���/9ݏ�k��K��1ia����E'&��r����cu�V�M��N�q�}�ɺ��G[�B��W�V(��c0�i�G��$�q��t�,]�C�������&R�f�6ko���괞���y�����7��lNO5@wR�a.��V�[h�*�����f&ś�Qݨ�dLWL#Q����!�N�B��]Oz�jGd�B�Hi����g6�"W���Bm�Q��$��s���=ٕM/G�7�Ox���a��RtΔ鍸Y�vqT��v�IX��j��F���s2�C)�K��W�X��5-ɦ��_L�6����([��Mp��f<[}.[��Z���T1��	i�u@�ͽ�I瞺��,JR+�J�4�{c�Ϊ;�����km�{�ӳ���s�b����!�R ƻEЃ�4�b�Ŕ*k�}����e�-F.����e������Vٝ �1j�?,D�9RTz
�QԔ}샥�g2�'�����XF$���bLA(�	'\�)U��J�ukwOX��7����I$!B�eR�%�ˤ��b�4\�D�8h�W4�����q���*@9-J����C^�j-�ޭK,���~0�i���@�p�\Q���^m�ALd���P��M��n\eL�5!#�yw��jBx��*��Ul&���m��f�^�'2�4�@�j�uuJ��۳��8%���J��.)^�Z��1����pZ�{��W��p��]�����2C��)���hY�T�]�&fp�ň9��l�J�=غ%س.���Z|*���NU<�ڝм���_�Zf�qjϔb��k\�B���sZK��4:K/���R꣰*��P'��:��O;���=,�O��	g��=��z��ޭ�M�t�M�o�B4E�f� ��5��y<�q~�#���97N�=#ri�g#�N>8�q�m�`qK�� A���j�7��c��΍�R�c�l�n�Q�o�n<}q��;A���t������"0�f*���ϯȏ ��ȏ&��8�G�x�����m�c�|��ۇ�S{��k'�>}$F�f�L��K�	�߮m�L��{{q�A�tGSuc�S�=�7ն�&��f{��v��|y��s3:�>�#"[c�.ft�#�\>�ֶ$=X�L��G��&�P�b�i��^�~�g�5�<M�|��m�巎�>�z��g��Lv��\v�Ht�8��C 4�*���`�`��5���|Oov�-�Gv���o�ǷgI�#||q�!�˛8��9��Q~�)O��T��@p��8�jC�l����ro�������q6����3�z��{x���\�;{�Y5�!�B�͢<玟&H�O�&�9�ɾM����=LrH#?_~~|��U4^>���V�+\�{��j��y7vr���8j�7{�^YGw��s2ep�+"�*'����E�v(P,!C��*���`*�%^�C�AU�-l�Z*�G�s��$ �w���ޥܘt:�a�*�YX��Tu�wBg-��f�1-���UBU0�0�!VLdROj�|2�D����H�M���ק�i#��=&�t�SAշ�7�џ���Y|�a�!���f'�r=���i�A�1�U�#��� k3q{7^|����G33��\c�;#�ަ�p�O���<��m�|�^�8�ä�K&| g�;}Y�\}Ox �F���oS8�ȓ��f��'�zM��g�9�G������~��Z�����25��&:G�q�� �n�o�8�.;��nCh��*`��8��ާ��*'C3@�&CY#�zp���ߋ��oO\��;uͤC��(h��GxžO��>M��sSq�����M�=\-���7�n�Lq=�!���@��!�#�~x6ae�q���~=8gH<��gDu7Sm����n'���۸��N�$3�8|!�La�w~Gދ�ʄyf4	�b�|�3�����Ř��G��f���~�����{[7���㷿W{z�}��a�: ���b�fh�V[gi�������X��@M'fh��5������S��8F߮��T;�Wה&�µ�ul�}��u3�ہ.���ibՑZ���*���T��#��( �41��4_!�OS[��t��Gj��Z��q��]ݜ�J��;��`]��5�d�c+ns�����6�C$�"�&�JGq���$��=o*x4�&�,qm�;��y7�No�n-�#~>9��=ysgӮ��!�@� �f�^^�˽W�D3G�ۜ�#�S�ӌ{Go^�c��z��{x���v�!h��}��鍛����c��9�7�����t�x�G!�>��<G�9$�&�:\9	4A�Ǐ�O������d"D�����6�}GxzMN��z����a�����q<B�38�f���W�",`s�(C4 ��ݸ~���{��c��p����#�8��ۉ竌~f��7w˓�GU�P � R8P�o�8��8�wgǧ<p�3�&|F�<���:~��M�735��9n����7�0��N�P�>��n>'��&{s����3���;p�M�7�޼��}����������t��ě��'{M����?!�?Q��A�!�a�7ſޑ��<EM�����i��|���#zz�zNN��n#O8�q�l�!��ā���o�~���wL<̜B(@�Ɓ� �7�=��q=�q6�$|�#�7�$�#�.�����a�^�W6�e.���/:*��!R�3�U�U�ED��tk�9�s=r�%՞�/��h�#�%�jK��i���q^��^�j�r��΋2h`r��Z���X�Cd�G:�!��f�e��R��Cv���4��_�m���"$Ր��:e�\���x��8`�S�@B=��x����gn㿴�qۇ�ޑ�D���t'�oN�9�?{u׵>���E	��FI�������zM���J���:�4C�'���~������� ��I�@�qC�h�J$��I�9��m�z�a^�x��G�� �HPx��C��8
nq}�6���{8�� r�AE�
�d�!'I�@�2'[��zv��F�Y$;	ϸ��A	a'�9��QF�w�zaU���4�>$N@�s�!Ic�A%I��f���N�r���%�"��p�Z�h���'I�5L���=QUZ���e���,���$G�q#��-�8�8�=�B��d�O�<a��F�T�<x���l�D��]k�w�P�A��j�ݼ?��\������+�S�o���R/e��[ivvV������,��E��tD��������\���=���7Z�b�2�^�xgG�d�{���,>��U�z�e6�3��r����KE�n�+d��~�"+�d(
�,t�d�0R���Pp�sG���,�Ip8�46i%i�0�_þ����͑A��G
r`q9'�YG�i��}̇���X-#c�օ,"�Q��aJ��f3�0�dv�S�q�9� �ĄI�E�"iAF��Ga1��������\�(��(B4r�H;���.-�`΋�}�9�7�Z9x�#�9���&����
$�D�O��7�˗������F� ��!A�#��)�x�@�iE�s3x�>Ǚ���q_�>�(RQ�8�L���,����h8�`����/���2�d!%Ğ(p���$�\�Nf5݈_z7�3�"S�e�EX�IR@G�I�c�+����v��W�ʏ�Oئ���F�t�􎁗��b7�����P�V�V3l5R�r��'�'�G�� ��Ǖ�Z�A'm�8A���d�;��&�>��-��*�i�=N5�t��� �%�*�g��<]�v�}v(~?(�_"A� �g���wlª~�i!�!B�ʵ$�A��'�$��9�̳����z8��H�r��'��9n8��s4�c:h�uE��T�Y!;QR�Ieȗ��	�p�G����V���T#Lq�����%�����J4�	����wI'��/�>-Ɂ���ҋ(��ʵ��0���<P����.y��@dIG|aJ��4�Ls��Fm����b\8���!x��4���<H�"�s��.�l�Qꉏ0W���ÖP�|9R��$ҋ��q�'D�rG8b�ks���f�aÎz����I�8�p��g"��W6�zv�w�`��8�HPx��C��>$P>YF�9x���V����3�;[y0<6�勳�鮖�Q����p����ɍ�n���l�)C���0�7sf��U☓PA�<8Ab�,`҂D!D`���ǻ�-=�N�W$�yuǖ)��;�)��:�+x����� �czb_M�M�w�{}̼�"���`C���D� (���=���j��� 0~ �,�����N{M(��+�:Bo|;!,�*$��$�J�� ����4�}���
���G�9Th�Q%�|A%Iq&�d���0q������F$9'Y��V��(2I��c�S��X����(Լ�^�i��O��q#��-���g�8��$��-�ިT��6�ׂO��.9��I�r�9��K��x�kU�mnr�q�(�I�8�47�$�M0�|( ��RA#�0i'�ߢߢ�$�k��)�-��Q�U� /�I�	̃�7���d��O�o��I4�Ba�J���Q&9p8�y�/>�߷���a!�Ą9��@8���	�[�!��x�G,�����f~�a�AWR�~G{�<a▿$��z©���<�Ƴ��F��T��M�<��ɑ.˾ɻ���t�ޡ����I���a36D��o���ӵ��ݴ�đ��ˮ���w���	+דFյԵptD[���D:kS��D�����z4"��5�#�"0�a�Q��8��cֻ^�����I�xr�H;�%�\[�I?	H�P�4q���ta)��b�'����Lq�K���,в||ARB��k�]a��*Y�L$�p㔇9�#I�J,�H�P@Q~%��֯q����#�8�YY�9#�����]���c���
>o�͍D�Pთd�)Ts�H�n98#���Xl=��jh��><9��$wĜQ�9�9-)|H�90||u}�~�΢��q�zd1�)�	��"�(�>�Qt���ب��3F��(�ϐ����Ƙ`�`�EHS�'Lo�i�%�q��q�2i�X��9�qe
���m����3�v��ۤ�a�߅]�H$p.H��cu�r_�gЊ��gp'~�{��O���E]}9i;�w���O=wJ�pݾ\��Jh����yVK$X!����&hG�k��}�\�o/wvU�NĹsiF䙽�#N��'`�٭ش�o��T��ziٌ�i�VZu�Ǵ�k���"4�T��	("�D6߱0ߕiC(� �=f"@z0kj� ������0!�j�I0�9�8���N"��N��0E �TDq�E���	�HD�Y��fZ[�E��W�*�$vn8�Fwh�!9�GX�ɿo\��|��I,��9n9$��#�9B��&��8c��߽_LEL���P珜q�=epY��xqʤ��9Hs�i9��k�o`%#�D�,��> r�AE�
�d�K�h4On����5C��x����$v�ҋ��A��Q���o��%}��3a��$�J��Gq�q��!Qc�3Q�Խa�Ǌ�3�0� srZR �#�p��Pst���+)�'2|QF��8�9��P�@�ÕD���H�O|��c�{�=���Z�oB��w��#�	`�7���c���M�*�oƒ�'�#)?s��P#����0p��=�����O[��=�k�K�z�mm�ٳ8e�|����MJe�Ӓ��R7P�v��nnv�k��w ��>ÑB�,��!�$�M*|H�h�|I&��T�'����#�����CF� B0v��)��J��7|?���&>�|Y�9B��%�s��e
��� �oqW��U��|��o�D�>8�D{�A�b�	)Ɂ�������g��s�j��97� ��Z�=��P��D�x��$ G34u�~~�*g�8�K�AG�(��A3�I�E�8�iAF�i��J�;��� v�C#s��e�FL�qG ��������8��9#�!�ri@}&�aD���^?�;�����>�(��$sG�HPi#��)�k������r���<Y�^( &��(����q�=Ys0}�?z�ɶ�ViF�|;	����A��Q��ͻ1�A�:�}4:ԞJ�K�[�
�BNN������e*j�I$�6{��OA�RF�\Or�ԯ7��4�v�-3Hn�Rʗ��y|z���t��ܖ��3�gWuO$����`�=�ohh�F��k3]�Iܽr�s�	�*r'l:�6\
��F�̻���5������1�[�B3)�K��]�5΂����׷s���Me����))�Џ}t3}|�U��m�;����N�r��-��b��ݭ{�/�CwT�Qb$��՗��=*�I3g6�@eP���緱 ��f��GM���W�aOqp`!�sZ[QF���c��M�x�Ƹ$�\V2�O�
���m+,#ܻ,���k��pU��7���D��Ը�Q�.�|���j��J�V��:&�V��uw�j�y0�B�p:ی���6�zT��Z)��1JC-�k���6s{�Zj[��L�<���uq��過W����-�Y+lJ�ش��IGɂԦ;8�	�����]��N�F�jF*1A��^JU��XS�k�p�X|㴾V�X3v�Zso����oӆ�)�خ�W�Y�Ǵ��W	�<�������W�����*�VT.�I^\Ŧ���ܔq��>W�s��:ތoh�.��z���
�R��Jy�#�����n�Ye˗���$�s��^I~���_��$������K/���[r�˒I$�Ym��/�����I/ן������tv�����m�II/��� v�wAﻺ_�\�09� ��Ђ ��p`��@H���b]�$�	$���r��I\e���˱�yLx�]b�78#�ف(!.IqrU|"w��2��{��`�YJ��OA�2����j��n�kյp�4��-�D3��oF�O3����ؾ,�Ý���D_2�;�.鍘�b�ҷ�(��zQ�DV����h����NJ���e+�5R�N�۰Www#�
�Suu�p��{�s���j!L-���X�%P�c�\��S�P���3�����P�խgB�ܣ�j[J�R�\`D��z��T�]T��ǉP�HK'��γDʇ9gw9�"B�����2+j��/9�������}H�xƶ�1��8�q�^�Qnj��͙j,S6���ǻd3k[�+o[P���`�����J���ڕ2M���Ӛ�*�Ur�d<�.�K2�=�M�b�@�˓�K��j,nr����BS�o4Q�{\�����;SL��e�M	jyh�U�	�� �s�&�@�D�]/2��ǸwW&�F�Bc�g��;p>�W��Eu�u �����͝"Ϧ�p-oE�$�g,e��}�sm9EA}��uY�M3�P�2�	K���;kf���\�o D�O�k_5���沗b��$��W��8�v�f���%��l�n�	�	/�Ԑ5ǸG�Ar.�m2�<����kJ�#�k�0Cr�G[�L`���5J霠��R����$����-�k[�]�I���+ڬ���1q�^#mͱw��ٵJ���4O!O��5F��:$5��r��
���Ʈ��"��#���t��o<5W
�	+nrn�H���#���ʫ.��sp�j��J�ލ�tJ��Ѣ�V\�ƝŠM7o[2��t&j����6�
�;����U�펂�u�M�#�Lt�QS�)������=��JîI-�-bvj#S�r��C���!�U�Y��-��Xe�0�<���u�r'«�0u��ѻA\�M���K�E��LQ���N�u�[��]�%uG���k�U�Ҥmko��~��6��b�BX�j֐��p�t�2e�ǡ�th�%Vܺ��+J����Z��u�Z�r�S��.���\˱�ҢK鑧�b�U�e���7�ȣ5T�u��Yl��d#]Tf����U�-�2���^�X'3h�Y�����:����~C�Z�)���D���kw٘\�c����4Ab�.(AYA�#���^�"sn��i|2��_P}5g=�:�=T�{(�Rz�s���_ �G#�����k� �$��I�ZE��y���e��P$�c}]�;��`���\�Gq�q��,B(��0�J�8b,�K�����q�<dk�KJD$r�@���A�L�Q'}W�눤��Q�\p�|X����ʢDt�$r���|V������ﮀ�q�4��F�T�<x���l�a'aŞ�&R<$	#�0C�8���e
K��!��Ĕx�f<r;[��3E��G�H
r`q���G�P�Ú5�S��v��fii�&H����8�9�8�=��iA0�
�@�G3L�>5?���mCA��A3��� q҂�>�Ha�|}[����j��59�qb,�0reH;�'�.-�a����׃����ZfI�s<�� �C�94�2O[aD�����#�>��}ՏԻ�dG	Ыq)��('��}�t_R=+kf0a��M8_I�F-_?z�,~d]1�qu�F��ϐ�B���%A�l7M�Es��3Uoo�>[��\R5𽦷X�3*�өwss��B���g��A(_]��{�w�R����W�E"}��a�>>d"I�P>"��>1Ww^oJ�_��i�χ�H��
C��<�%��E�p���'�����q����_�Q%��9�$�F� s��
�ak���:��NWQ�;!!��I�F�]�@�P��N������;�y��5Ϡp���"�,s$� #�$Ҍ��f>'.-k���b��`�%�H(�rU�&���8�Lq�sY���qD=��OI����ʢDA�Ahr�q�q�6����Ϲ����c�I"���S��I�dK�@�#�#�!����3�uP�Fb�ÎS�Pf�P��B�Q�L$G�
8�녪x��3x�<@yɁ�������r�I}��Q�5�q�������f}* �Y%P@�AT��c������\}r�˩���i-�nE�.�eF�xB���3��*��Q�ݶ湬��bl9}��P��Љ�*�n�4!kS���4��5٫.:Ɏs��w�J�����yM�a���DX�o+�:�:s��_Hm���y��M�����/"�h/M��$@ �*�:�Z][��s��UYw�G���Ꝓt��ϊ+a�ގ`t3	bA��B$�E�8�iAD�|I"�s�=ʾK�MRK�L$!������ɕ ��&�\[�H��B$�Y�f��������|��q�r�@d�m�c�K��YE�9�6Q4�=��+ѝ �P��?ĐR�A�"[Ɣ^���P@s�g�o�ѿ)тh�A��z%�$s8���0������^%��y��3J1��46�|Q� ��
U�$�E��WvU�NN�(-�[�c����K�	*H�iF@�8��|f_uz���k�ܖ�D�i��"�A4P}$��1�)�	�,EQ���(����|9C����H-[�!���x��`sQ���O�3�k��I�ȗ���P�0A���Ӊ�| T�~�ҭx�p��n%�e�θ���{���}�;e�U��'�ݓ5jj;�ƈ�(,�]�c����:d+
}�ݮ�����sLT��
﷦l�Ԫ�S��(�Xx�ё��7|���v^h>'V�NVq�jV�:�+u̸�����,(�rW]u�jnN[�Fb�c��ޯc�0+<h��!zIGǌ$G�
,��H��1T@�l�}~G��3H�S�[#J,�χ*Ԑ�aBs �b��O�H�$0̄|9�@�0��P<Ǌ$�.O0�g����.����ù�V޽�t���ӈ�˧�^>�;�Cc���"�8
��^�~�g�Zd�"�>� �D�(����S�� �|8�YP�t[3Ҭ>�2�$��'�Ig�H�ÎU$(8	3��)�~��a��i�r�q8�o�(�%��P@M�(��f.}������Onc�x�YY�H�'>�J.�ds09p?Ѱ���A--d�Q��d)T|�8"܈9�k��%y:}19�$��4�J�>�O�21�$����G(�� �El(�u�2�G��h����B~]ѥt�\�$M�4NDb�Ñ�w�C���oM�cqt4�Ah���c]4Q��< �q����n��8٬N:��T�RyQ�e�m���V�Gi�ܮA���p�����wk�/_ �� ����	/qOS�n�B���ʵ�9{�[G�/V��w����~�0`��r\p߼X����s�}Y�]ֻǂ4q�Ďr�CC9�<YBc��K��I�4w�B�<x�ȧ��($r�9��K��w�.Mfk(�s�O���1���CSu�QfH�|( ��RA#�909��pxž^������!|H�M) =�aBs qA��s1c���<Q�iR�x#�H)ʁ�>HD�Y�4Wr!9�M�ئ ��
Ɗ�# 5�q��P�9�6}d��﷩W{��%�����k�"(���'h�8�%��[ϜF8��Ė`Y��p�BH�!� �^^�˽V�q8�n$�J�V���=�IC����N��.���U���k�s)iX=�ނ�zz�WV�+��ɍ���YÔ=�2���Q$E(��ؼ��#Т����s-dX�B�hK��`�Hv�C����SO��qy���"�)𜳃�F�AN�
=�u^T}��@�re�!iq� �.�C��t�	'�r�Y�g���ɝ�}�P�܁i�I�����}/�<������K oi�;	�x��vBkCa#��|>a_���SSLH@@�$H4XpA#�-ȁ��w�D�9��`��d��9��I���JIA��Q��V��X	<���;���s����5"���!�
�t�H�F���[���q�|�hg+�YBc��K�<iC�9�������\ǡϊ�����9.6��\��A�ś�>�R��<�şa����A�b�	)Ɂ�ru!A�6o����w)���j ��$��L(Nd"�4��4r�aV�E��S{ƀL;1HS2~$"M(�M((���r��"1�� v. �;,���ȕ �ĚQ�0��l:���n6�sa�}i$��V��BU�A8�;g�`��6%Ȏ�9]�˫윱�v���#X41��'p��b�C�{r��T��)wF�:k]^a׃mS�1�Z���Q:V��	�ǲ,�F#G[�:����h����ENU��&f�vhL�#Ɇo"� Ō�t���g�7�,s�"+䜁�P�lAn9�=���z�z����D�8,�G<8�Ѕ��9N8�\�Kiq}�6ß5�Y*�Wy�$��r`rN�I,���D�y��N�ڈ��Y#�;	ϸ�
vq1�����3��aD���Ω��o���Kr	nD��,EX�QR@G����~��K�A�9n9$��9G@��C��d���._�誊����q���P�@�9TI�Z���=g�}
�z��hg*K<YBc��K��I�dK�A�s�px�i�9b��%Ƹ;	.K��!��I<Y�s�-��ul����G
r`q9>HD�P�O�o�'��W���/�z֬;h�P�,ͅ����#��Bǁf4�۸���]5tV�q�����0�@�>mϺ��U,�CGMl�&N��p�p��\�I�]6�Wo=䌓quVԿJ&9���D��y0���C��t��C���$"�` lݙ;/[W^	|P�� ��6$r���0�h�x#�3�x���診8��^RI|Qd �PQ:�8#��#6 �u���<Ye� F�D�qE���36t�n�z���ڬ�I �I���>��$��rp�q'3t��K�}|���0��rhB�	�9N8��-���Y�7��:b~�xl/��9D�9�LI�8���0�� ����P|���In�!47x���d)Tk�H�0�j7��,V�E�y�@���,EX�(� #�$Ҍ��;���΋O=G�>I(,��0rU� ���I-�%����q�r�:8��H�qʠ�<P��q�4,Ұ4�UU\}S�Ul_�^W �~p�Ys�P������Л��w�ތ�nz�U����C�c�]�yY�qO�,!#�
7~��X��uv��}£�	�ԫ=�V�!��݆(3�/F������ʁ�76�m�I�-'��I:CЀi@cJ|�Q�>��vk����Yc�!;8I8����.9�9Bጏ��o�b��H4�ϫ�.���!����,�	0s�9���ԒJP� �p�&#$�D�P�*�	��<>��8)��v�K$qϠ�G(��,s�D�$���dIfx�^��� ��$�<Qd �PQ8�8"�G_�}*<��|WY�Ŗ GÑ*A��O\[�I�S�� ��ks���k����(	���I-�!��Y�f9�I|��l��{�h������9N8���$�J�V���b��{�_T���Oi&�yɁ�:�,�����q���p�7�K��!�5qG]�@�Q�H��r7�QQ(���F?׿�S{I�ٙT���r���넋��֫v��9�J���q���5��M�y��3�v�0A!�	���C��օV^d[[ÏWl%�^ǎ���I�{}ٛ݈]}�U���7b��4��r$%ƌәD�e*�'sי�Jh1�n;���p��n�Q@���E9��T��Q�9�9'`�o�=E�y�)%9g� EZ�	��2d�Kq�q�ۥ���9��R�X�����4q��2N(r���qGX�p4X�I�S4��ω����DcX	(s�ϵ�Ez�;ks�pA�2z��ω>,�9��U�H$p�m$�d\t*���Q�8�%�$��4�iI�w� ��s�m��>�=/3���$��0r�	�B�INT ��l�=Q��z���s�đf9�"iAD�H��q�23�ie�s1�e:�>�*��8#�ʥ Qp9n9'�S�� �I��a�}�Jt���O�tIn98o��c�,`�!(X�Bo������l�+U��ɲ����ex�U�)u�:��Z���M:͜Ќʕ��7��g�W��e@\�w��twX�a�[Xk͑�{��Ϟ�����t���ws��9icw�ب/#(c8��9l^�c��g.P���5�*[�{S�vM"H8V��+S�y���(��O=���9�>*�ծ��a���E�-��_UpˁdS}ޯ7s6m�0~��e���!�.��]R5iZǷ���'�>=]�x�e���ӹݯ�Bb}/LV:+�]��\b4�B�u����Kf���bJ�^�>se�IJ�Oxl�ܠ������a����v����|�7�&Z&�i���N��6�K�ή�5��湃'�wa�=�WZ\*z�[���{�,����l�a�t�-��|W3&gh�=�̧5ڢKN�� `<���{�gC�u2q����1��N�"0poe��x�p���,�J�.�_R�2��Яa�:�]Cٔ��{	���`��4Md謻��U+��u�P\W׋��f����'�����u�d5r�ӡD\\#��|kkER�����e�Ƙ�]��e����{��;��:v��xet,����ǘ����b)݈b���������җ��]X�v��d�R�۷�[$�K��Av��nݻv�I$��%�IrI.\�rI$�I$�I%���}}m��}�����n� ���������� ���Yf`��{��}y�f�����@�K��%����ym���I$�����!( ����<grbz��\:�uT������nη��t�ڛ�_�<��{��D<K,QN+����^Nɛ�G�b鲰<���>V������F�u.qk0`m�(7*fN�a1�5��WES72n�ǜI�V�9���8T��C��#k���\&�j�]���j7�M�6ɡ����cX�͋i]j���Oo���!}H�I��oP}m�Lڤ(��緦)�mp�鏕(2���sj�Qdy��k��C�o%�6���P�b�fq;ЊK+�v`�:w$�ϓ�>o6�]�ܗ_m��eZ0(��ɱ@ܬ��̼֩V��2*�lJ���n��hqх>X0u3�w�#Pt�dd`�G��Y7F��Ɋ�%zp��#ID�`�7����O����z�Z�H�\�|1OP;���L�{X��ů�õ�t�*��ɵ��+OC��0���MY���9q[;��a�S}��k�u�.e�ظ_,o��Nt�����D�!J6uV&�c:�.�.��^8���w�/�a�w��N�ۙi'd&x,
�}����Ƞ�͊�V��%i��^�T��a�z�%�D:'�HT��*\T���GN[N�7]Tfh��ޚc�4qBi�i��w��W�u#|�j�XI:v��E�W�����,ю��v�M�6��fP"j�H�6�mL�F2�����2��J�(��O�2e6C3j������=䝇��ugv
���<v��"�QP���ؠuQ%ʾU�*qtg�7�
���_\]b�f\�?-��ÃP�P�2鐍H�Tv�m"g!C��T��էH�#�$8^-T�/E�v;t��yۮc�U2�W��7��7�	Q�*��� +i$ht�R�����{ӻ«0���²�*��D�/���븯W=����AlZ�\P����s/�YF/أ�U,�)ʎaT�@�%Ij��P]���\&m�y`�@�NU�(��kuە��XcD���F�8��U]R�I[oܬ=���ؕL�zԆȑ���t���ԛ�ں&�L�q�%!��	�c%0Y�`�Cm6C4ᗖ�q��������lGcV>��"���!���#x��R�K�U��s-V�"ŜiRN�D�~�RU�ȝ�rfln�����Ch+���+�g�j�Juׁ�l�șr���#m�A�Ζ��îF�rhè��U\���cx\�u���T���n�)r���J]��l��]�{�b�&�Z��&�*��ܭO|�#�$�7(��HN�7Ŕ��ޟ������6k���J�V@���r�(s���Яq������=c�TIdd@��s�$����k>W}
3�65aF]�@�Q�A#�-ȁ��w3Xl>("�x�|xs�(��8� srII(>$r���>>:��?nWzˮ��B����I��ᛥ���,�χ�oQv����3�Ĝ9��CC9�(�eE�C����9��7մ𒇏�E2<�d�P�@��l}ė<��-��v��}y�����gĘN�=b�	p���k �<a���J�+rRH�<9�M)!�_qD�<;�}���6E���\A�&���H�*M�RI|S�!�9Xp�fv}���F���Rf�ɶ���_ro+*�87y3�2ڂ�W׊�Y�:��Y��`�@b�T�9[1��,�c��`A��癋�K��~A�E�l����e9/^񦈜*^/v�����������9��S=6K���ݥ��իG�� �P�KŦ�@$Z�I��'��f��Wx��a-XL���Ye X9�]�=c�&��m?%�琉+�=��9�$�0V�� �,	����g���R�������G�q�@�&�F$�߽�u���qQ{D�����B���#`}�{w�?k��U@���H�G�.�'�I"��	����J�o�(ߏ�J�����A
U�&[��qb(��H�F�x�>��P�|Q�d�<����Lp�!U�fj�R��?�}?^9��lX�Q����XahAU �~*�5����|���A�q���XQ�eX�M$���Jv\7=bp��XK��.7��$���cR7�@���p��k�\)�h�n���VDc�m��}�ڽfI�F����i��Wn�$:�x��8p!��g�D!D`A�h��c���x��\�,��G����CE�ޥ��S>;�j+8�(&䨏Wa>�r���nE���oS��n��$�a�'�\b���ue����4�<I��@�U�<O0:>�IG�{�wu\^w�I��(��ǂqϼLh�X�OeBߟ����f���$S�&�RI|S�!�4��4���Jt颏��t6�q�e��`�J�w�!�p3�)�O�Woas�tu~���VlS�"0�| wZ;��p��lq��X�Q"�Ҟ���������zR�4���� �P��F��d����m�U�B�HO�T���������3=���T��;�dW>�b"�Ivs1�'�C�D7�I:%H�6*ǲdC��F�^Mf�1�k}����W�U��;ef9}ԯa2`�0�}��D�
yetV>�m2����?�p��.��F�fl�r��v�O�|\�AZ��%i\��c4��AOh���\�V���\*�
<�;�R��*x�e5�r,�&��\ڲ�՘
LO�>���&�"hV)��#���2�{�g��,���8!V��|��4�A�s1�%�|{�I�<�B���"ԉ��4�4����Q���5����
P��(�B�%w�3�Eg�����-k����q#�#J4�0x����bd��g���8]�IO�i=����ߥ�<�?Qœb�%C;��iR�j9����v<�i��6�}�PM*'+�=�M��0ʮ}_GuAS_;E�������[
�*��
0ɂz2�;Q�c�M�Pw�Q�d`��׆�}��ha�9����U5pQU�/5$V�s�sGC����*�C��<����-��p��3*tb���6���_Bf�8��V��\��)�nLHMJ>Yˌ�6���sH;zP:����s���]��v�S��&R�3�-�|�a��g9�{wcu��"�X[�ϝ!uh�N��>&�Ov=K\�9����{�{ٓǱ���/�&��I���u��y�1g����0��(WD��DJ<3ch���ua'�6-�}�����|�msٝ�w���/8��Ji&��M)Pg���Q����g��9�M�D��jD��ƓF�F�����A1�>���T�I$=bO������b�8߾����O�f	P$m�E�$��<=.a���=��=�&��I#��X�I课&iØ �)�/�3B_33����/�h�J4X�|�n�k��s�U�p--���qщc\����ED����ǹuA�7���R�&�7
��V�!��߄P#�	'��y��[4ht%�]�X�[����o"�!~�Oo׽p\ٙ��YΨ�M�@��^�*�xq�րd�|K-`C��2�;;��ݬ����z�\�ƺN_���}�t��(Ы0�Fӫ�g��)_0 P��B��)�A��o䨚N��a�l��}�a�4��O�(/���d`�R����S��L�X?8sCi�5��z&�90+�j��������h͋��X��a��i6�A�}�^�黚��)#M0��4}Q҄��(B'���8����Te��x���|�G��kG�[�<L|Ŧ�e9dҕ�E"�)&Cc@>�Y�n��,�o>�0�����d`����xz�2ŗ���h���Q$�XJp�}>�ɵ�w��ق��D䩌#27��sq��f�5X7��l]�� yL\�>���r��좂��U�s٘�cD �ph�b�/����1�ݵ:�4�En��ت������KP�T�H=ۗ�r���P'�*�.���0��{�fȫ���2i6��9r��՝v?480pv0'��Q���}����r�g�2*��IN�"�Ŋ��ᏺid����tu<���Q��p�h�Ѓ炸�>т��簨���=�M�x���X(�H�
3�L+���w_A�""{Eq4%�&r+���[�ܳk��6<	@�'�G�~r:�w�b)c��q<|=��M/��������J�t�b<8zŤ��q�ڵ	G�GI6��]Z��n��>���@��6�ࠚ�7՚��]����+EjH����Э4���;��1��a	 �׿l��R��q�[��T���R��[.3u��T�S��uR�FC�Jg���B6�o��P�Y)WN-�8�Ȯ���(m�+���<�Ő����G9�;�Q����B���OV�5�+�v��4YD6$��%�6]D+PCĝ��DP�+�I2�#�(���=>z}�*zԉ�.�"�,�
I�9)�p�G-o��� ����I�S����N$f��34u���Ċ��D�f��tI!
Cw�	��B�_E^Q>���W�L
ӆ���ɱa��`�~��6���,V�26�?KɑT�������%��\O�Zm�(��
$B�<S��B����������*&������څ��^���[|�[����,<F�Igx��hl4�i��+d�!��.�!4��P�%�q�ٶi�
0F�r��ִ�ȧ�#6�ӈ�̘h=�H莅���X��Od�ө�j�<ىvf�ϗux\�kSG
(V��m�7ysΕו�ԫC��%]�S&14l�ۙR�q�8���u/r�ǻck�����u4��Yk���f�^��x.\�1t�Da�]EJC9�k��g�<M�q�H�G��]�瑻�Gt<z�j͈�>P���A4,�t�Zs�����[�Z�����.�i����M. ������\�_�`�+�dg�&ԉ�0�n����(�h����I4'#�T�I$Gfϵ�ޮ�QS3)vbv�oÒ[���<Q�Y��[��t:O�"�DE�JSgJIOŏ4��f(�,���� R��YV,"T3�OA��>�B�޻�1:�%	��(&�9�"�0]���z�z���O�
�|(��� �Ѭö{b�B�m۬.ͅP��װ`���­�=���� C�q����Q�1*�Cß�n9���^����<�����(PP�B0EU�!��Е%��Ŏ�,�r;�R��NX�<Z&�ڝO)8�tZ{iZ5'�̠w-���h*�����G绗�WVj|��u<���+�x�$j���;�/I�(�}@V�����ѡ�"u����o_�c������T����c��ͅ�lwoۓQ��V+r`U�Q�6,$�g� kg��I,`n,*q��"�tM�4;칎碪*��I��
	��!��h�pI�>����ffr�CԖx���q9�iJ�t�fl$��E��7�z�� �=�ڑ2Fi�(ә�X/tL��g��'#
yP.�$���c����܈No�~ۯ$c���#J4�0x���Әo���E���C��?b�Ig������bWw���<���C��n4���Ν'��#"��*)�{��*���8*��>���Y�qGӻ�֥׏>Zc��QH6��m�\�k�.�OV��^�v��RP燒;�!~�d���>�d�y9�!�\0�j����.��	M�*g4!��WpZ�0��	dc��ܧ��8�w�9�\Q�ެ��}�fu�$��u2/�{�W2��y�kJ���oX� �ǐ��Gh�1����r���Ƭ[����֮��=C���o��m��_st^۝wfhY�={��q��Y��J˦����8�^�îvF����ޭ	��J�~s�Y}D��r9X!�E�Rz��;s޾�����j�Õ�\b��}v��1���!����'��n���{�]у9*W�XH������]�
TH�쾚����%���ݮߔD#�阳F?����*�l��{���:�Lk������fb	|�\f��̔�,�k�FH��H�6�75����Owo�j�K�(��vad��)�H�@���1F{he�n^z\/eUˣt��3�/]�-��L��D׼�*�Us3J7������ܓ�*<��j�͙C��-U�k�I�fF��iࣆ���kZ�-ʘ��X[���/Y�
�RV)��(ch� C/����$�9�?_��I$��JK������d���������I$��m�^��m�I%����\�r]�w_Y�����͗.K�%��}�ٙ�>������m���{��s���}���/~��nݻ$�ߥ�}ق� �I ��U�0�Z|l��E����.�������e�3�9[*P!�UU���ZXMu1��s���ٌ�N�[�l�ӝWQ���i����ի���WqE--���"TOPD��:�,����}ڷ,�EX%��=�1e��S���M�jY�Gk��e�wR�i��Q9r��ms{hf櫥���db<��*_Yf%fij�[�C*&rbfo}�8:�����&�޲�({kB�6����VL}Δĥ�b�}\�ӥ�+l"�MQ��Z��_k<���5l�o5���i�aJ~U�.[��L&��ՕA���-��]���v�(�8U)	���%b6F\F7��b��SFWqzq�Z��k�tn���vݬ�C�i�i��FgnW�)R��r���h�O��ĳ��z�S��E��qu�/zq�Ŋ�V>���g�έ<ЊJ��V5���.���Gf�f�]f�;�Wţ�f��I;!m�uYA�q�QE�{��)�EԻ[�ۢ�@gJ	�Y�p�z7s�L�n�Q�
�}�f���+��|���ŕ]h=��ܺ��n��;��V�1�+�����Yl�I�qn�ۣWFZ{��a��tu�7�_)D����¶�U�-�	^	&Eb�eT_?J� �˪^ȃJ4N�?J#e�gUڥ�^Dzl�yIS&Bu����AV��]3�W�Ĺ��6W^�j��Ct8�̯!��u����8����������R
�hN����l�5�ӷݱS��8p�h&;'��3e�z���Tv�q�H�Aa����iN�J�!Z��;��\��A�.'��Q?Kmb�� [i�]����]� ��U�q�x��oJH�D�dާ=�=9��x���sCf�lȉ�ʃ�k3+�6J.�Q��R9x_��}��a�ÑF�c�)Y�B���u���j��G�:�V�hʪ}YR�{Ņ���s���F�ea�y]�B�쫥��!}��Y@�0������
�xu����6L���Z�	Y}�}�Lj�ևk��TS ��q?r���A�Q�ꡇg$kwȣ�8Y�k�f.���	��.=3LR˨��3@�ۆ�о;&sH`h��M��ѐS���yr�{R�����?+�i:�U��cD( �hc]4h&�C��
�Ia���e�j˩F��Cws]�lJ�Y�7��3n��A�Ӌu�]~��=�O�i{ȏ6�;�n[lJ���mYՕ�y1�yq�(��Y:YeX�D�gM*\���������SP{Ġ�TD��"Ӧ�q���9r�{o�����D�XE�����-�jU�>΋'��~N�|�&�(=�Q�0\�9�t�ޚ���d���;���M'K�z&��0sf�{9g���8��ž�b"Ť��N�Q��Wp�c��u��{#⏈�]FT@��Xj�>��,�	�	ɐ���� N�i��I�\�n묹�,���i9dҕ�E"�)�cꞪ{�^��K�Ln/���~$w�C���wΧ�7ӯ�l�%�Gu��uU�"�7�����Ŧ먧4z��*o�;���̅ˠ�F��M�V����x��SE�A���K�,���շIt������֗�tsT���t*�t,S�3�5N׸��;�CbH ˪��it79^����G�������>� �τ!5�
>1"�P�"4<�$�qMx�HhY��0��"D��AC$NO�yP[�$���<Jv���O3}%�n�q�~�Ɖ��P�e���5�Y�0�����4_�$x�,y��Vx����k�#�����'E����<M*PsHF��c[���S��9�_5�Ӧ��GX�`�9�����=b^"�zPc�[�jU"���,��o^�j�["����:���'���͹~qį��&�z8�,z-�_92��4���d�̬�Q���x8
&��4��x9����a%v�Ѵe�&"�tMT@��7��A7ԧ︺-l�#���o������`?�g΢�½�+n�<�p�e�usV�i2fi(-�uQ8."�4�媮�q�Q�{���n�v�M"Z�\{z��oaq/qd�.����B�[r5��x�ӆbk���;x���8�2��'��䮭]s��N��e=��w��Ȇ���Pd��v9@�@��X�1X������%��n�^0�R��C��JI��hÔm����Y� �)$_�Gő��hNG���I�r����b�j�B��Nퟸ!���ɟ/[�W�H�#�>"χ�T<F�JS{y�4ϲ�7z6�粒EG��(�k�H8`�Æ
���X����˷|*��M*P|��jPk���.�ϗ���i�o��B�X(�H�
8�}�ޞ�+�D�(<��_%R*M��N�5�����Vr8���Ef�B�0��ٚ>Gޗ#��@����u~B�D���q��&�P6�mvӷzf�b�.�=������zQo�#��=��b
���xp��ޮI ���h���N+>����;�4��(��;N4�e��m�#"�q:D�;�w4Ց����2%/2=e�	����H��(&��@�&�eD?&�x,�<=�M/90*��Ϻp���s�yA5N8,�Ty~�?
`,�c��������xe��0��fO��(&�Ns�IgG�^"~oHvY\+R@��iG��Zi'S�����<q�^PfC��JI�؟����}�{9g׬.$n�FF�I�9K��mi�ٱ"�<[�RH|�ħoO�9%���#N��-����8<ʡ�8zR�>'���f�Ŕ���}r���R�߉qZp��M,�������������8肋�4�x�&EY�����ګ�d�j��lEgQ�� �J��ʘP���Dir�o���=��L�wJ�� LV>˓�\�F�K{&I0���(���Ǽx����ڤ_9�[��Yy���Z��k\��շ�D���jF�	*0'�Wl�!�5[M�'��`зFBQ��ڠ�=]	ѣ:� _��<(�}:�4*ł��G�~fi9��k�o0�4���_%R*M��Y4�k3�{���?MEW334�IxC���K'�t�P&�|4�`>,�~>�+��3ŏ�D��&P�s�ň�Ğ��/]'|a�C�ϸ����taQ�,WF���Z�ѿ����}?��I���(M�ࠜ,rd>�+O�T\wϱ\����((N�aG�X�4��s�����/|�&,f�GQ"�)&C���L��T�fr��os^a�N#���`�����x<�B��y��wu\_Γ�i�����tg�iF�e��+�nW-2NdTIY���@n2#�*��5��FM�Ѕ��Gi�ܘ�G7/Ş]����=�
�1��0!w�6�a
�88p����x\����D�x���XV�w�Ws�j�h�ӵ5.:o�uSi��؃��*V�oa&Xb_pkt�0Ъ"���72�En�|���?{��j��7�Q��ВG��X�I��8�r�iTD�3��/'{�&ł�N;��y��>�O�v����+妴�i_%*��_!�p�n��'�딼�3���L
�h�D/�=' ��c+W�Ռ^���EI�yM(P{���?1�Q��[�F��xf0���O���M�>N�=1�i�ey���~����M1k�X!���ϼ�'�О">`%� �F�G�X���� }f'����ɛNSϙ�U���(&�����Z��w~�����`�w7Ɵb��O��&��7H�3]r�~2H~뉱j�㋼�UQ�(7r��x+��xP�,S�O��pU���%��G�&�)���VU"�m	=[�n_l�������v�r'�o+\)����]�з�qg:m7�v`<���Y��j��-6�=�T�$PZ�_L�,Rf��GPE�V�8n\���#De%$�lM��L��4�4�c�Q�k�x���P��K����!�}a������/��F=�v��In:3Hҍ"�eP�p5Qͳ��ޖљ����R�E���M*2��|}]��Q`��K���ɱ`�S��x�T�&f�����z����u�������J$UFEyI�gi�0�y[�wL<��>�!Q��A��W�p��a��| X�7zф҅|G!���f���HZ����30C'��)@���|N�=�M-r`�a�Tb͏�ѽ���`�>�{�b"�I�g�tҍy�^ozk���/�V��.Z�$���>��>�b���_��.U��fC�������ܙ�����!��]�nR�'z� ���t{��TH�u�R�nE�-�gk.=ӑ�|���7�F������ǮL�tc�&�
T#�P/!
>-Z�L�y��"=��z	�>.f��$Q|E��>���B���	�zy�c\��:`��}\W�jH��pȻ^�g_�y�/84��R�I��JT�(q�O��V�}��</�EF��jD���(���s0O}p�A���>�����B��<Jv��DOQ'�ޟ=9	�����#�,�<<ʡ�<=.a��_ϧ�����{�I#ġ�(���l�	Ƒ-�X% >��Q�l\&�Ix�iRrg# ��l�s��/�f�I�[g�_!�:l�X��p͔JU����W�5�/���d"<Ey)"�l(�#�铑
��/��(�����uл�33d��8��#���S��([SW}�sҕ
ˉ[�{�%�x��0&�|9�˔}��#�:*�ډU�ZX�$)�W�3\��on�����ɸ��b�M��%N5���(����a2�>�-[�rn�:뜺Jw�_g-�CD�|-�$������8>,�_��
��]8?�ިLߣ�K��Bnti�6X�[�4�ɁV�]ٛ�9X���fc��a���I�g����p1��wW��n�`�����]D�E(M�Р�a�0�L}.�f$�Ϥ:��� ws<Q��Z���ߗ��nS�a���,nA+	�@#��򡋸�?=�� 8�(�?-�&ϋ#$М�9Se��;����P�*���I�S��\"K�7ľ}#�0�	�I�f$�E)M��b�߾݈=�����͘�>#��U~)�I�op���Z��2�Y��N�՝���B��S���5s����KӖ.�����H���:�$�4rr�^G,W�-^�����6�� ��jIDC�M�Rm�m8t݊	��IƲ��ڬz)m�tQr����-uyr-�ڪ�m��:�(��V`ӗ���N��@$zȢ�E��Rc�0���D�9d@��,��z��~��
��L1����a^J$\3|afC��lC��I�g|qb*����f(�_����u��Cʂ����%$Rl�"��j��v{�f�|8PZ'���_D*�is����K�M�8�>�z&��L
��]�9�>�W��LG�x��Ry%���0�Ԑ$ai4��~�=���W�ĉ��'"�	���c�7���Z��>4'x�� ws�x���u9�34?�B�y%�|کaTE"�)&A�{���q�g�N��+���dEAA��a�0J��G�"}'�z��n�eU����5�e^���nI5ɽ�xe}9X;�Fevթ��[Z���CUns�WP0�J�n��u�� ��W6�e@D:5Oi�1���e1o��Q	QR��"�ϢE]2-ۈ>ͳ�ncn9}R5�LY�}�{;�;���e{�C�v�a�*¢V��A�T TeC6�e˓~���{H�n�3K�Q锚�{�[�ɧ��E�٩�˲+�=�a(��k�z�US1ev�H���O4�{��Cj�ko�O�zo��d���v[���7����n���Lq�n�S���x�0V��S~E9�߷���Vh�Ƭ�]Y���Y���b��q�;��n'D�*�n�Gt�l�=��*Oe�Wѫ��b�+��0
AZw;�Ž��k��iR��Ηb$M_:\p�U�X�{�#6��y���%�F]W\}C(к5�OR��] ج���)b�����k`�\�rŒ�s�;A�*���f����Sc�N��spCymq��M�9V�0���'�N]9k_��{+H�N�Uݽ�S��~��F�٤���
�}R��M����}w�鼨�p�R�2M	Ų��X�P��%S�pg����9M	[j�����G��̺3SR�,p��@��f���ƕTת��T�:
���K�C�!�uf�6�n�K���nݶ�I+�n�l�I/���۷m�v���$�O䤒I%˗%˗��$�I$�I-��6��/od��v�۷��� ���������������{�G9�?~wwG�9����7wt {r���엲Koo��l@ �e�5�����[�Ô �Z������+et}x�7ޒ�S���
�x�ъ�ߴq ����}֩��H�ɽ���{*��K�4,hT�ج�[�Xۙ�=��<�:���Q}��㾪���Ыɯ���,ު3�W �%�[(�Ω2�t$o�wQ�b�L+6U��]���Vo��
f�B�r����C[F�绒�*�:�iq�C]�P��Ѩ�W�tP�CfK��*G���uqu&�)�@U�
���WK_'Ƚ��Գy:_t�|V�Jsp�RV�\-5��B��p�=��ո�	XMɞ�4���N�0���j�zӭ��������o]kv"4px��rŹY}�²����p/�������П&��C����.��i�VKk��GV��.N�z�]������9��m�aN[�5�b�(sTn������V!�3Q�hW)	�r}�j�<���Y��Mlf��A����ϡ��v�QEJ�t	�TgJ
��gHF��-�[�Ű��B���P�Xz��i�۬�P���OF	�^+1H+��sC��l�-�;Q�nB�fB�eC�w�?3�#�f+@YD"�!mU��W�X=�Ҷ�����9?>HݲA���4ޡ���7g�o��{'��ńk���GȾ&Ö�oS7.��Q���h���A㩛l�RZ�P���,�k_��7:Jd&1FϬR/���3q�U��$;��AWp۶��ݤ�=LHI&����d����3V`�J�""q��w��-��(��	�wW�����Q��*�;B�Ha�{���m�S'���+�d�}%�ᙞ�\t�^����8И�wE�����C�rE�(��̕v�\���"��B������(Ca4U� �$�6�%��94ڎ��f ��"�u���:�Ȣ�7n`�9F�@��H�۰r"p��F�7�YN�G#~,��.�����Ք꩐�RR��k-�d�cSC�BP�R�G'sی�R���`�`�y���=��#�}��U8,!�`��cvd���]%ZY�6� ��#p�Ŏ0V�t���úz�O�����7���&�wS�n��{�	}�Hb3VN:u���\���9]>�U�P���i�S��Y��^s��@�ڥ�G��d��S�<�՝^y�N�康S���մ�=su;��(�Gs�z�Іt%`�����̱��O�����-�Fi~#�w�}�9��ࠜz}��$�E�����Bs~�ݱL �Xh�� y�p�V,s}e���ު~�$�2�)A3�⼔H����p7�>%���'�ح6�M�v
H�H���e?���1s�$~�|EZTE&���&�-��\�ӟg�ex|�160p��LM��4p�|��]Z���>��b��&J �w��?33�X���-�|��6qE� H�<Q�,WF�3�F���^�ы�" �&�`PN92ZWOFw�(�/d`P:<;���ბ+G+�t���w Eͻ����:.��ί	�[�<qA�V�y���U�4��B��$,��Ye��HA+	ת�0��6�/�r�ϸJ��V�I��l�E�K8��bz�fUl�_DAP�0tڼE�Ƿ�{�+P@E�gH��I'ޥ�>�׮x�ۗwr�u�⮬rSV���Gw%u�]:��[�n�H%0�:#2�g�[�0־4N�x�
�Zi'��K�.��'~�0_�`�+�d6>�"�	�3Q��ߧ�t�u��H���I4'#�T�}�~fl���=ܦjg�*��17�^%8��#�E��j��Һ'��i �Ľ�J\v�h4��ET{Y�<*JzmL�3z�qJp��8�lX&�Iq:W0|#��]�]|�	aF3��Z�H��������]���z�z�I���|9�
H��'G���[S����a=j_I�qM(Pw���?09:�w�ӷ��1���2O�R�6:0��,{3)�_����v�r="`�ZW�F����X�u���"⒊��5CwU�c�q;I�RzV��b��X/ɱ�Xa�X�h�4Q�����n\�foV�d9�IO4ⵊĪ����Ĳ��vs��j�Y�2lVV�xK�K��B��]��G��� �IV�4 �O7�AH�	5�9y1i�K�h�w!x�$� 0R������{J!4[��`�xJ�/.��������f>�)IE��E��=Q�\�s�U_ �M�PPN�92\V��Y'����8a�r��T�x���q9�iJ�t�	$<bԾ_0�ǋz��!�ՄZ�2Fi�(Ӂ�Y�����|03@�^/D�|*���!X������<��ep0�&ߦ�IN:7�>(�,(��}9��$��}�Q~ jX��Ad�cȪ���qs�o��Ql3yHk�Y;�p�Ix�(���dn�z���<��Al�`�&h���f��8W�����ٻ��_�{;��1�ܼ,��� �9'�x�u�u�ߡ�*�%5��~(���O/+ �c���Q,7t_ٓ�����]�M�Ι�w.���w���4�Yn�tE'3z�Q@�vn��"A� �]�FՕ؅��2@%D�-Q�XD�IH)%"c�2I	���U�f�s��a��XTXc[CV�����(����5�ɲ�M(P{��b�'��k���W����<���"�	�Ѧ���e�K\�9��Q���護� �����b"�'�]���J9����v�<��r�D�#�X���* zP�F
�>��+c���l���u|W
Ԑ's4�$�]�u�\֍��M',�R��H��V%<1�O����lU�Uk!�Nq�L��<EY.fk��K��5@��˹G4�X�)���'�o�����Z˿���[�!��X��I߿[ݯH���g��e��T$��!��h��&;+����ȇ�>z�P�*\�����z��t(�������Х2&ꎶiٗȥ�|O+˝���7+8�����[���7T���TJ>�em������4�CG.���.֜����L@�^"����-�F)K�d�dJ
��P�0f��_�;B��1�`��5C/� h��K���G����q���%%�>(��#f1�z�+�¿���I�gx�lr�'�������~���/�J2!�Z�I��ev�V��N��A�e���`�xJ�x��Gso������q8X�[�6T
�l����q޹7sw��a���"s�Iv�M(�$������z�����KGº*�� zP��ࠞ�RŢ�b�4���3���'s8���sU%�ݺJ��mM��'<M)Pg���V%0)s����}u5?As�옴ȳ��0�o\k��wx���P�����Qbwjb`K�7�3���L����mVrRҽ�ō�@� c���y%�*���h魓�Z��>�i�r�w8��D5v:����8�Kz�&'�Q�"Vd������sv�sjܑ [oqJ�fĜ�wҳ�����@�"��(���QE�����r�����!���_�����
��=�g��qU�h6H㏈�|QE�T㷷��>�n7_�U:Q`�*��JqRp��M,�f>��ױ��M�xc��RK	��PA���M
�����vL�����q&���QE�Cx}$�E��6��?( �C�"�J��ޟ�d�0Y���:���mP�����=�<���� �f��p��$M΍,�<=��M.r`T�Gi�7���u��O$�K��IJ�0�0O�و7�F�?i=SV*��V^0�蝻�Z���y�f�N�ŷ���h�������R�k<����*�W�<7�X�h��H���DVۨĒ{7w�� z�vSF���a�����ɀ��$6s"�f����nEƮ������q �2M�JC�0PSkr�������o���Bl�
	��8�*��������:I��'s�Q�X�4��sI�*{7�!%1+��a8���.l}\G�!��~{�p�#�!6�<P��O+���h�O�gD�Fdx��H�Ğ	v���$��i���ȶ��� ��X�QD?���4�dw�|���y�����|��+��� ��id�	Æ.����������Ii�R�r�Z�Ъ�Ej80����⏙���i�8��	"D/>X	9��|��M=�>�i4d�,J,��臼x�P�Si��J��Ȯ�#g�#6��4�ֶ�nڠ��7�=ȲEj���v���9������(��Nh��c�i$0y��Y}�9����j��w�(�vޑҳW+��h!�%��Ӎ�u 曗�АQ.4����n�ޖ����;Dܖ[R����%�V�@��N���V��>�c�O��Y>N�T���I�(�~>�+��?�=K�(���,D^$�3YEh�O<Fx�g�6�-AG�q��b�8a~�_�7g���G�c�*"��6炂p�ɐ���?�D\wϱ=gG�Y��	ܬ(����~Nx�Z��^�dL[R�βQ%jS�>��j�FoqD�g'���5��8�>>#E"4����i��Z��~�W|0|�?ŻWբ$��Q�Y��=_5��x=����D�sh�,*��f���j�(�>��p׾0�s���|Wۦ��wu�I�";�c��x�q�^uٛf>��?�O�W�p6��9�e9=�FNC��4��2��3�G-�U
�p���=n)R��݇���p����gz��N�JNu��}O�d
M�ٍ��Yk#t���o�r"����u�HL�\�(Z���{V�[X���N��>�J�08Z&����g�}��ؚp�a�6�N�Y��"���lG�y���l4JXE&��Y4�A�#K��Q��[�U�Uy�`���Y?O��Ό4�,{9��;Oy���z������\�(���,D^$�K��3l���'��fi��( H�>>,���G;��4�]��93iʘ��*�_����;�o�����}�޽뻮fa�񃻛��b�ޢ�x�R��t�f�0��޹��fcÙIL
\}��m@�#<ih�3|j7���x|�m,x,���S�?�i"�'�4�m�:&N�c0@��1=o�fX�&N�g�*������ �<���[�g�!=�M�{�_�\]{���/U�� _+����י�RH$�[c�=Ye��N�5H+�Jd��"1gs.o�:^�hژ�=\i,�k����}�5t/6��s��~��])������`15F�"Jq�~#�"��*��$6��z[Xf	G�v��N=
���\�����Qc0�u�YY�p�Iq>(��3QƩ�W�~�u�� ����ѺN R):l�4����Ի�	�01�a$@A��E�20:�{��b���b���FT<�X���f���HZ����1�3��T����:X�[�4�Ƀ�j|Y����{�u�ǖh��"o�<���izQ�6u���V�a�AbE��E��z��r)Bo0{�D�+��.C��0x��~�;����IU	�ꅗ9�4U���7�I����!}��[��7��]l�pr	Ǳ��Z�@Ү���|�]˅ ��v���p�3�X���b�2��y�[�ǢL9�2�;k$����]�zzkCi�Hg�p���F�=:#�dM�����W9dYq)P��)G|�ؾ��m$�{�5%U��+M�O�d�D�LY��X��k�ϗh��'��)U)�G/��/�b� ]<U�iU*��Ƚ|����C���N0v�>p�i���7U����nt�ؗ2f�KS��"cb���|�0j����zם	�on�="�¯Nv��r�f�s`���<�k���!��2S����-�u\{�k6�Nui �t򗾰�T��8��,&S~����~�ͼ���W2���ڤ˜�^b�IY�(���E8���7^�Kp��w��	����6;w#:�L<sgtD��WL�̝j��_m^�V�����[���o"V^�J�1*�W.�-�n�iڋ�x�hY�/'G2���pP����\	�_.~�ȮI�޷��ؽER�J��m�����9"�WW)5��˾���+O��5���]�G:nf�Gw+�`ٲ�uVE�N1��4fIR���Jp2)Uz�[s�̹��4�)��\�X`��]��ʢ�ۺ�^��\-]�][��%,js��mڻ��A����P�4�I$�I�9��K�K�/$�JJ_�om��%��}l�I.I$�Km��e���$��9�������~�30Y��[d�I}��kl����y������s��9� {�����Y�ݻv��'�Ѧ�݉$��U
��uRx�D�Hgz�H�
�;�Տ�e^i��$��+.UCx���+�mc�n?����3`��;:�q�n��Z�ًc�����tS��t�#�(;��ͤ����+��tH0n�I��D}}p�(��*Zג���t���j�n��I�Z�����\��{l��7nF_19���\��5���T�c��J���$b32.wg$�+f��_)C����yS(Z5#}�`=��P2�Nc�]����b���]�It�Bݲ�r����M�������%L�Le�W�GWm]��EDN�v��B��mf."w_}��H{���ꍬ�X��3Y�/5:�/^5����G�t�a�R��z_��R�*�wm5�}ut7�f���1�Xz�_&�b�����m�a�k�5TӮ(Uz(�Zŏ��湚r̾V�P��픺��2�K�¯RW"d�	"?�w.<E\��h�R:�t��E���ᵨK�u)f*j'v�lKK���	(�%,�<��}��w+٩>�[n�.��I���:M`�j)��������B�����wi{yi,�Rr�NA���ig/,���8�pUY|��ѨH_J�%��S�j<z�AUI��NQ2?-���̅�d�T�z5kD��%�)�5�4�<�cd�=�DR�xY$.x2�XB��Fb�룧lCH�ٔ�:�n)V������4��r4U"Ev�0�I"/P�I�����6�K��$�ͦ2��6k(7t+Ud#ec]#�ot.�Æ �e`�-ā�@�܅DO�!��9�vz��m6�\��C:�C�'嵪��D虔�V�ɉ�̓�����ꈮ�x�z��k%�h����f��P^:�Y='o���!7W�B� ���AR��NHj:0�-�2gf�gtaJa�}͖	�oS�]<"��wvO�K��(����f���:�#Us��d��%[JV�[v.��ҏk��(ŉ8Id*��ي�j���̈mba���%M�T�&�x���\䪞�T8Am8p!�ľ!���hѧ�&��cUݻ]�N�Ϊ����ъ�Yw���*�3�cY[�`�oLy�,Uj,�1 ��qx�َV��yy�{��5QB4�R����+����V�}��</3
\x��m@�#�E>`��`��!j�1�<H���)����Ԟ	v��DO0�I���O����F�QdY�袡?���$����<3^���8X�*����'�A�Ty�>wX6�|V��"R^'�)A�a�|z6������t��?��"���q���O0}e%~����_0}���X�����+�Q�xf�Ӭ��k��i9�+�z,�`PO%�*xj��혗���v�F���e�K�T�fe{�'�z.����(י~�:�&O*�<�޿���MeǊ��i�k;\tuWf6Uo>���/T�(0�.��I#a3=�88pe�c��G�eJ��V2jI.�f��*�f����i<��[(��/K���^K黺�����Nic�#×L{.1Ixi��Gl�*XΥ��K��K��h��h"/�K��ҋP@�f��OuO���湛�ǬQ��=bC҄�{t ��9��FIlI��_9�M����;��b�#ۿ.[Q�L��"ɥ)�>�Q%bS�6=�z��j�o{����2Ex��>0OE"4��b�.�ߥρ�Tt�zĞIv߫�I\3Q�%��"0���(È���!��%�ol�Y�?n�2z{�3�a��`�
���N*N���O0L|j�y�^%�f��ڒ�|QJ<�9�y)�k�E��]l
��Z�����lr�$�	���y^�{��t};�f�VM�_%�:��cú�~r���u�9~[k�4���+'���.�o��4b�!�7O[���I���ťsX�9[��SU�z��m勋u���|�6����}A�������g6M�H{H&b�E��Ax6j��S��fI�UD}��q��=w<1�,1CC�&���E�? )���s�~��o[�}�qbχ�Y?�T�#��6����G���oD��ɁR�:=�0!���N�TGǈ�O$�?�^Z��#�K#�,�L���~�~hiQz$=(L����p��\�y��ծ�>'��j���U�p١#I�>�]�$��j��D�G�J�2:�F��A����N��+�3��ID����=P��O+���ŭ���I��!�Ry%����tf��c��쇄�p�A��(��#D�a9�1�j��}�eEX��hA�=z�W�-�t][5�U�P�z�˝�.�6~`����wU׬ON@0A@�,$�OI꦳3��$kK�ƭ��xb3!J�]��,Ag���Nm�M{*v`/��D뾽�U������$�����:��f���:�ݷ"������<��kmH�~�u�p*��<���3�,�Tv�M\q�$�}E��܇>+�M
�حG {��h���Z��<Y69f�D�^"x~�)��f���]}��:!ψ�J��ޟ�d��{�/��_Is�����,��v�'� ���V�jiP�t1V\
�l̇��E�O�3�X��Ih_!��P@��|x�,WGGI���G�ݕx$}�&s���p��R紛ә��u����y�Xh����
�NM	&ְ�Ԏ���e����%$K�Wi��~�r�?Q����ߏ��r���.�#����9��b*�6�Sit+*�w��z��YWɽT�P��W}VX��F�|a&Ig������
�q�+�_m muELS�t���WEK�}�d��C)�X��`�r}J��noj���Xpe�\�r��D�;X��{�պ�3�ݽ��7vn^���A�8�)�;���ȴ1����E">)�9�dC�͛[��ǻ��T�RO�;}u�S���4�H�ዽ���t�!x��%8����X�*���%=tL�z�qJp��8�s���t���}�B���g2_|�9�)�UEyK�����!��2��ɯ��|9gđ"�iOI�6#�(�������R��Mӈ�J���G!�������~ɍ0È�w��AN;c���ǳ���_�sٵ1s;�k%�J �Ӝx'�J�sͳ�'B>��J�E�~�t5݂E;؎�8R�aj�/Ə��}xe�Ҭ_��չ&�{�
G��k9�&�	�*��I���pQ�:��3֨��HX��̃Y0`��8*��S�L��:�6� WU�H{�ŷ�!�R��яoޭ��e,�8�Z�A(��<ŵ���j�����r�ɼ������ghC��@4��Qḱ�3����M��A���R�i7�����>�����;�%�*�8eRH�6�9�2p>Z���B�K�K�XE��2�&������R�}4��O)�2="�'�FoF��Ǟ��16�4"Jqѿ�G����!�����FE��E��bqP"��ǡU�ᛈ�b�Q�מ,�w���<QK�k��ݏu>eM�x�r�q)�U��I�g��y��&�%����ᤒM$���)�9�a�s1�ﺥJt�5ɮ�$�x>�<X������d��Q�~VG�Mғ���n�Wof
K�:�K��*\�:���"2�o{���j}}���=�Q�U�V�����x@�����LȚMÍuv����U������fi{�ݯ������m�&]EΥ�T.�cpʲ��TҾj_^T�Un�	�y#�<5�j�5t�[�[+|�-�Y߾P3�t���6g��>����C��AN;k�M'K�z6�"\�b�Gvv?�v߸o/�As�z'�J�/J8������r�D�#��ȻOF=ؑpBm���w\����	���������<$���0Y�]���_Yu]��'
�IM�NA��#�X�37�	No�諺��؜�-4	���4h�cьs��	�����S�\t�zĞIv���͇��zz�^]�}�>(�,�袈3Ifx��ގ��Ed�8X�*�/�8���%�w���΃�&�N),'�����0�7�}���i�-�~}nZ3���M�CW�i�m5:�1J����{�S��p���)��A���� |�I
$�X����º.�֛���o$���9t���zP�\�q��3ob9q���20vI}[�r��Y��@� �Y��n-�nF�>Y�����f�v��F�S=A�8���ӡ_�_��n��Egp�KY���ǥ����s�������&����=��ݵ����p֘gY<
�,�giQ����{`��a�賉�Ǳ]U�S��	�}���
j*��q�v	�R��KҋP@���E�k���:C%a�
3#$I�{�<��E�ŚX�
��&�{O	!>p�qV��	.�/N�Ӫ��I�S�g��ǬJH�=���r�sj���$�jh*�	���Ǣ�S�3qG����"_�ŝ"�'�]���E>�'7�0i�ۋu�F��͚��O'w6Er�T�/�g�┳�R�uKU��	)Uq]h����mw	��( �41��4_!���n�Mb���x-��ཋ�fn�8���-T�wJ��ou�T*K͎80�^nԾ�y���}���r}�N���6���9(S�[�n���9nG&:��u�z��Y�b�[d&�!(^V�LR`��2b�iz�*������g��E�T�G��R�^�����E�� n�� ـ6+�|��Lr�X��aH0�%bӐ|�9�jSBћ���2�����I�o�x��	�K>��35�p��o�]��.NY�i�TE&���I�5�������o��A<M��K"Y��*
�bτU��|�7:4�l��+���)�r ���pf����P���e�e���aV�8c��=޹ߕM���$\��� D�cȸf�I���LLDO�ޓ����<$�ix�RT�+�e��gg�,�1t�={�s�s��'\�i�h�v)ey޺�j>��]��U�>�*l>�e+����Nݿc]�Gѡ��Z��|��X���발rgNo/v]--�ul�ʮZ�Vh� :,�#�#���X�#���\W0ܑ@�X�ad��_V��!-3��վ_m�u���u[�Ě����|�:��Y�W��}���]U4�'<f#�V��.?��'����s�o�Y�����*���ŋK��6�0��$^G���">ĞIv߫�II�4�8"�~N�ŏE	��%3�s����X>-e%��S��~a�a;�T�ݦ�V`�8f�8z��O������Iig�Rrr�Z�Ъ��j#��>>�������_	���lr�&E,�#�>�IͿ{\�xx�	^4B>"�J����k$�x5�5ۿy󟦪k��cǨ��ő,�4�)�mta����Fd�9��0W$���e�D�nDG}��yz#䌸�������L<3�\k����H��#�) V{�k��Ww�/�uC����"�,b��!�sr�E����ݬE���T�mb��L�6��9��݊�Md��UK�}{�]�KVR7�jg�8�����+] '8V����v����ܾx�u�ɦU�q-��^�3ً;nA���ߪ��o�kyy�Ԁ�(��)��:#P3:�v$INY1�q;���d��gz�Cw1w�W�hт�������VT���^��鸂�jQ�ݕ�B&��YӇ�h�4�؈y�R7D��ĩ)�\�8��q�;}Fꢼzj���> �T�M�o����kpsVʼ*Sٟ|�Z6��1����J�V���w��w�Gf҅-�jb}6͚��]tI��y���Dڮ�2d�����"��I��<���k9�}�,[���FB#�!
�
�ŧT,'m�C,k��.6�����Te�ܗF�Q>��<��x}Z���!n�r�d�
Zp�7ф���'��V�jmu��ֲ��\�/ ���C��㎸v��#]_sY��:j11t�͆\��S�F��X���ZyI�x�n�����ߍU,<��:ׇv���OR,����'ܨ����So�Fv��*ˣy�s�����;��۶[m�n�m��$��v��$��wt�v������$�N_��I/�\����$�I$�Im������Ͼ�۷n��wt w��ww@����������Y� �����s��ﻺ �}��h �˗�6���/d����m��Yy$�^�����/<�|sof����_U��y�5IZ�SI���άꉥ����+|�aK�,�I�N�;�wX-l޸�bObs��Ior�û� �T7�Xi@R���]]���T�TV��[UƻvE+V'i+�yw^�IU)�u8JW�Evګ{G"L�hᰭ�U;ruC�c��Kz�ܬ��[����7�������r(,�ٴ�!���\J�^v>P"�e�:t��O;)�c�onѝ�\��l<K ����=X�ᆯ��T��鄍���n]���g�����+e��R͍���M�i��c9�1ݬtn[N�#�����v���[lv�}��r�U��8�h���B�M5�V�QJ���U ^�5]o^o�w���hR5oz����x�v�آ��I�U�劵WJG��3��M�FV�X8s���˙1�ͽ���<19�dZaS�V�j�>vIYq*8��6�[О)��/:]QL�%��6�Z۾o��}��Be�!� ���/(Q}r�}�����;�2�V�u���;���En�w�mA�Eo"W�N8:���g<���U;A�Jv�U'V���Ʒ�\(�'����Xq_�Sk�Zr�KD��dY�%��S)Y�4��tA�O"�)�ѕ˨�! ����h+�'%����oY��2)�1�ʖ%�vFEcL��~��@�G1��]�%׆�Y��P�gQJ�xeH�'e?u�^�v�mm�T�zAI�j܋kº��T�b��P�tDݯ\E^|�9ikW�r�݆��ii��@պ���p��!9N��(qh�ƫ�l++���.�uh$�0a�뛾\}t��WuSُV����B ��m,.t��.�xG1�,[am&��� J��M�CK�h������+3[g.�D���M.��e�e�&f�q�Ķ�,�	�c��' �$u��n�b߃��Q%�R�e��=��CcM��%�U�0�{.���5l���,�H�����(Qf�&�jUl�N�&�<�Ůߕ&I1Ro)�&B� �KU���i�0&�r�&ǇNH�q_i[I��glaȢ1�B�ĺ�$�_��M�t��]��Gv���6�9v'r��s�q�+��:�^`A���'V��=���ұ4Y�x�vϝ�����}�Ь�W����nY�-1J1*��'�S[���(�G���U�33h���,���iZ(�OB�?e���߲{慄�+D��Bg6��cȥϸ���s��WY���`�T��z�(���>�I&��|��,����u�#�Z��.?�^&�@�f�{�+f~޳������oE"<S�r��"5�ּ����P�����[�}Z"JN�Q�Y���k_j�G��#+A����h��UGp���\�(P�������YY�p�Ii⫘h8��w�{��s88t	���5`݈v��>�}�v)׮R�3����"�"�,�#JzN@�"n:����[��ׁt�������5H]�t�i�Q.M�9!���i	fA�u��B��C��A�ƌ�ۿ6�JY���Ml�t�yӺQ�A#;Vξ�dI(����ޠ�U��T\�A(+���eR��D!�Vo=/�� }I0O��"���)y@�JQ�S(uBg�F"* \�`�Ia�6�ɥ
=��.�0��-��r�@���9���RS��:0�kRz��d8{_+s�� ��H�ȑ9��	�M/�sb�b�;�|ÞO	!iYi��.4��3zrf��Lx-5�K�Y)s�&�{\�|]�wz���䐻t}>*ԇ��G��)�7I����0�z�R��,���sb눴�&Y�I�G��F���<>[�g�G������<��c=*��{����MQ�II��G�<E�=Q�3D6��ކ�&ri�i8X�*�/�qt��m���6���@eڙ�}="��!���'*V)�N)�1JS���{M���!wW�]����.�o����e��0XBC$PЌ4!X,�b��{�Q��+:���*��|��娗�ɢ]�oz��� H�̚�:.��KT➖(�!4��Q0A�H8���� m\H��0�C(%�F]�0�u,
}�K'0Oiǉ�K��xvguӱ�V d��DՃv6^}�M�v�W�U������񅑢�z#�=' �C�E|��d�d�=})���M(PA����쓆k���q���B��AVA���kR{��۴�s�.-s��=��do	������8Y��M�rO��Z��RB�0�ȫOG�v$\�����:�����9D�D�\���i�$'���.���Wy���3���RT�4�R���#�X� k}7�퍑�I��Gv�i�L��ѣُC�L*�~;��Iw�)M�Vf��Y��խTi�qj����[j
��m������F���-�Oݗh!����I!���v���˨���$s�"�H���Ņm����u�-�gY�wzWm�F���n�v8`<*Om���	UCh�E�D�z6�:lGޤ��	�*?R^������l�����@B��F�l��T{~����I���O����ҔQQdY�袈I�/��{�i5�|�>'��T}���4��f�G��Ė}�'�4���Ҥ�r�Y���0g��W0������g��l��iH��>��q���a�_BaE�6fl��@n��8�+���1���?�O����O�)����(���,?%��+	Wa�봉r��b��7����};�=������zYi�$.���S�ꪉF�&����v$\��v�K��Uy>��r};�dK�qiF<�����]f?���Db�,��(��`��j��h���"z��w�l6t�@�L-���A����k�lͬq�j�]o�����9J�a��틬y�h-<�2�#��5��Β.��~��c��✭l{�cM���l��Ϊ�4��D}m)�o�B����$���� ����o��xI	����O�܈~�7r�9��b�с!h�"��P:_���~�5�y����XCُE"4��.��'~�>|,����<��W�������I��x�0�,�䢈�*	L��a�c7rd�{�f�:��U�)
��<������]�c��?�mJ��y�s
�SBя��!�.��:+���M�w��0���s�g۞��G����LC�^J�Hg���Z�mg�{w��gCx��_\.E��*V����<�J��:r��W���i�zcNz�-�S�kl��gC��:����}]�+��ӽ(1��`�G���cnvR�'q�A�3b���fC�]:%��M��:�H�7z�qDz
�V��bQ�v��*��X���G���,��#��"�g)_�"�$B�/ȩ(��h��`�PQ���A𙤫��m�"!h6����!}�Z�W���]��M/����B�>4�9�6;�����J{�"���o� �0`�� �\���&!	�|�a�'�	���!�I#I�bb���y%�w�XATL=jRD���� �7��w�ySÉ�ID���y袄G�r`�j8��k��B���!�Ry%�:�%'�4�c��w�ٕ�O����DG�A)��8�����gw������'�}G��eIÞ�I�؛���,�Tw�&����Rrr��Jj�ѯ���u���U[�E��5r���f��{퓆����o(i�G���9F��A�rn
�Ƴ(&b���*�����\�IR��Ǝ hѢƎ�����4�*��k[I��"�f�X�%O��ט�`������$�#XYr�|�)X��.&�L�P�ˡRQ5D�)-!P�:�`����
b�Q��4�D(�J��)��n	>h�b�+�M�N�R,�)g�S�5L���Vզ�߄*�E&Mb5�j��f�^�������\�?@�4{%���R-��F�����UT�Q/��ZD�nDz{���~�����}Ec����qe�����4�*�ѯ��j;�����>�9�d�D�\��zp�f���zq<�,ԙ=|=U���G���]I�q�r��ŕ����%$K�WZ L���vE�O��w����(D|S���������犊���v���$��F�i`��b�53���#(:P�������qPw��qH�v7����b��
Z��"������H���._m1�$3,����,`�� n�6ް�c3Ҿ���ύ������L��soqjZ�P:Ր-ɕmk�r�HU#2fF�H�}CwEnZ���m�&�A��E�SK�4Q'�i#d:Uw�0$�(�T�mDy.h���aж!���,zQ�'�k0�|�g�L�y��x:�'�'�4���\3|Q��p�����|X�*ɕEP���g����}�}R��xvR,����F����G��b�jq?��I����Mdڅ�x�N;:}|�d�^+�S���h��=����Q�ݿ{6�.g@r&�%Ϝ� ��كؚ_�`p�6�jt#�m�JxI
�⇚O&=?�7f^l�\+��� �zd�\��K��ޏk����>��]��0}i2z���V�2�$x�R��t�+O֯޹�}B;N(E�ڂ��%��W��Y�ڮͭ�]"k�P2��7����xjW/b�ǽ�1~u��(h��6B����8y�ŕN�56�����B�Yf�wJzP]jÊ.;ҥm�R�ܝ��w��X�o.ҏ����R�"��e��l�,�F�I9�&R1�E��.
P�RP�PTZ���� �ʡ������KH�2=XAh�2�&�����O�0�m�7�<a|S�=�'�Y��Q��OmvW0|�~��JN��x{0{(�#Nfm �d\v���jF&ri�Y:X�*��'���qW�>��� 5�ON`���?�&�.*�w����s�1��aؔ�'�����q6A�4�fo����>�*���B�|"�z_H�=rO�����)��W������
>�|
��5���R������z�.
�g}4�Ԟ�z6�"\�Gvv?�v߸<��As�f�bi��,����gW�s!�����dK�ڙ����5U��{Xz�*��Ӕ�U3|k��䇚�6�V�,���Sx�`���IB4��U_��oڒ�X��"���z8S9M]w)ʃ3�'\�j�N�N��l��e�5�a%j��䲶��P�L�l��.�n�P1L"Z	y��V��!j����2P�Q1QZȤp�� Dl˸��8���l=,:��b�&�3]��zQ��Ð�"E.w��j!&w�#�0�������*h��pz�$Y6�A�L=pAr�o�誙�@����$�@�{OF�fIp�K�I=�X�[��"�'�]��[O0|h�v��^]�hz'��G���<T�d�gi���ɰ�G��ǪOFx�kq�gFCvKǢ(�8��=��|<M*\A#�p65V%�}qE.K�R�[E�d�B�f�8y���~��	��>zXA$Dx��k�������ez녲����s0��S��r�p%}d>�G3��y
��K�қ/������B�q�ǡK���KoK8Qj�३&�_��W�ѷ���Q�x'l����~�ڹi:�vy����l+s3�el�\Q��.6�.�z��;R-��-;#&�e�4^������Ӈ�(�e��\ڤs�s^Vɗ�u�˗�B'b�k���%Bd9[��	�?B��9Zy�C�.��R��X��T�N9�'��C��(�F���Ȕ��:���7����e�S�˰��N� ",Sz���5�vm��VCWI����uD��uZ�B�ۂR��F����P2�%���8^�9\륂t��`�7�K����c��Ս�3�����d^Zݒ"��	MѧJ�~��S���Q�,�>!����v�xL�H�q��ںb��V��{��O�Y��,�Y4��#m�32��������R��λ���IU4Yl�3���۸�mZ�RՖ��#f���,�{:�,�=��ܶ����)U��zP�y1�$�=M�K�[=��qo3�7*��Aw9�{ڳ��ޔnq�M�a���n����֣W�3��>�j�>��^���������i�x�b�B�t�'��Ѿ;�y��WH��*_e��Ǖ�Iq$]z�Βi0�,��$�ƒL�s���%�/�K�I%%/�nݶ�%��}l�\�yrI$��m��}v�-�I/<�)����s0�3m��쒂7wt`뻹�I'ﾒI��t�z��   �{��~��w�F ������A&���P 뢧��V�̪
��Vk�]���×8���c��ݑBUy�0����ˬ���g �d�"GH[���W34�w���;�W}�����u%�@�w	6�O=R`{s�;z�CL0a�U�f�h�3Nq�֣y-���Z����(E��V���v�C����ɍt�t�k\VP^�e�@gZǉ�)=a��eWLWՏ0�٬x�j�yI�!N�����p�LUi�{ܚ�.O�v#���٥gj%P��"W�o5#_�*oHz���q۸is�C�cNґ�v�m<9N�$�q���B���,8�-��*�����f���-ޅ7to{��7���[WWn4^E�S�k����)¯�ݔ���o��*�N�Ϟ��nU�
)�^]��f>�:2�sF]���3�Z����ʘz��r���j�9��^1��h����[d[�l�1���4SL���[�h4�gKf�7L�4�j���˰���/l���wvN9wj�';�nӭ�p���UXGTG80VL�Ζ�������Y���|��mIs���G )df�}�m�`��p�1R�8zq��P��0��4r��y#f������lZ#*ȉ E�@�a?$9��9(褨���k�M	L�X�˴�gR�l��D�uSf�7{d�L��H��dX"c����J����J��J(����F䄲��<K�*(n@M� �&���o��Zki4�0�^T����y����c�J ���\0��%�U�pᣡ�a
�-ڀ�w1�c����5@�j6Q	 ��o�Ԃ��w�Ն���3�N��J��73��%y%�e�0C#�DG��y9*څ�Dn5��i�eHI��:Q*�N�`l4�֤'3�98&�������#�QS1N��"ID/]��n�-�8�2%E	Vc��B	�&�/�4)�!<@�[�6
F��1ц�]z�����̙������uuȡ��a:Xx�u߶�"���a�+���E�к���I�e*aHn��^d(ԥWZ��e��=$J�9L"���]
�r1֩m��-�N�!a��*�]�օ�t�����9����ZؤKa�\�MQ)�A""����V����4A�01��4h�U��NvfdzU�޸
�*S�����*���PR�M�`���!���h���	����$AE��"�:��A��ۥ���b�JB�$�1Q
@���-y4�@���( IR	$O��P�1J��ԡ*�B�P�PQ�E�4�B�)�B�u�]u;�~��u	��d������Ϳg�I�g�3��MbOx"��$T�� W�m�z���ڱ��	���M/�������c
,{��/��o�7�OB˱"�ރ��9��z:�}����o��;�Gjy��ˤ��]��揾I�T_��ǣ	"\������l��<y'8�@�Ta_
̲(�Ҝḣ���?�1�T|A� �I�%���m% �c�Uǧ�z�*�7I4���>��(�*BP@}��RΞ^����B� +0,. Ʒdi�5�7��Vv\S]�K�j~�5�q!��g��z��yD0W!�a����v��0-�[f��Z��b�`�뽻�C���nM��[�J�.Q�yr��p�tTڃS�4�7P܉��Yܹ��,�b$0I�^{T���i^� e�\.�R$�'�]�d+�@BP�b���v�$�Jl�v���(��N�F�PHO�u���2Q�P@S�I���͵�Ĩy%P R�-���I�!�

E�)��$w µ(&���4�t}(t�h��h<�lq�"�,�Y�Na�¯������NF�aF�W�94�=�5�Z9��ݽ����i-'�,�,�q���+���E\-w�(pw��=�9v9G]�H�DA�Ә�,��#��y��P�%�
����XA��A�7��f{�{]�ĸ�{D�����ad#����K���ɣ���!d6O��B�
�mi'WMo��)�K��(�,��$��(�H%̓�.�>#_|����﯆� [�|"Ͳ
(��0T���7n#��"=�_`�5�m�8��<n�wT�{�3�z
��ZvS����� C�u	g�SШ�8`��A6H%UR��:��v��ŷз8���ȹw;;�nRV��D����R�N��Z��U�eV��k>���?,�w�����@���)	J�)8�T�S��H�S�!1S�4�j�f
��N(D)&Q��$	%a��JHAO!.��6h�(���\�J��E�1�Ʉ����ZNI.�[IH2i����ƜN��,r�*T��~K�ω>,s@�Ŕ���M����NY?k[���A�i&`���5��ڿ}>��~��>E#$w �Z�I�<��9��|}{�u���Q�E�Y����9�4��[�6?b���h��L=V����ίX���Xm�����k��8�F9d�s4�
�|4����2`���䜿�(˴������,�� ���֥�|o!덲���_q��U�(�8`��j߷�~�����?@B��rG>,�DK�q%���;���C��:o��8��g�>��Oy��QK��v��+D�ϫ�W�彸�S�=\�-�øF�ۥ�a���r$
0Pѡ���䖄��m��Crɝ4r%�5��.����_(���.)D{�,r����e9j�l��a����U�	��I���$|����I�BP�`F�I�h+�RDB��h�(F�IA'��
h$���$����Sl |I. �%N(@DHD��YU)�|Ì0A¥ok�sz��D�h((!�3$�>�Z9����xɘ��Q�Y$9F�A.}x�C�k3{�*6~���{��<Q#�
(��0A���k1�y[����_%�|8_�[Ih2�4��0s�'��o�G��<L
0����ğ94������r�j�!��v󃆹qd��r�>�$�fh8��O{��y��>4w ЋD՚�@�=��@|m�o2Ib�<YBf�A,� Ҝ�i�a���>��u�k���p̦�KD">�O4f�0�:ݎ�EV���>9����
G�;ᤕ�9v9y�ӳ}n�/eߢ��kS��Ulſ8=���}���&
�,��ۛ؄K���ʅgP+hp�<4A��pA_P��������m�� roDv�]��ֵٔMI�T:l�q�xi�
ʹ?=!C*�i[���ZH�2��m���E�ٰB,�>��AP���H�$�����"Jb>gŦ>�ϟ�l 	1��*D�ڌQ կT!ED0�%#"��I�Li(źj/"�D�j��S&"D�d�YcA
�_��f��f C��b�Y�� ��9�-|�R��>i���r- ���*Ӕs�bE��WvfoNLۺ��3���$r� ��|I|9h�o����^����&No� ­ABQ�-� �$��>,Ê=�K� �6�� Y�(�����S��g�4�)�`��}�Iȑ�f�-^F��=o|��|�b��M<9fYE@�Nf*Hm�Ͻ�A��S���X��r��ks�����a(�\���L�9b	�R)Gw�S�;�Ǚ���>��M)(�=l��i������Dm��P��yc��Y�n86���{�s4����V�2S�P������(s(��"_^�+j��N�T��h�t{�1BA@�[�����v�\��Β;�3k��V��b�\#����m0�u�R��k����wx2č��s9ӳ���u��Q>,*jHK��� �"��i ���B�Ix��mI�-��`�M�|	$�qѠ1��$��Y�BHn��$Z�@�"D�$
� I0��nU ��s�r���㜪��|䲸��v�m1'���ʃ)
#�&FW�9�|aF0OF\��6Z!t�p#�N�+��\}u�P����"�w��%jN]�Q�i9�������e������Y��%�Ҵ��l&�9'��-|�$B�+�Zr
>��.v�o���-���s��0�DK�q'�9hxI��'p����w��W�e:�DDIh�A�$��(Á������˨}(D�w���8�z�(�e�Q\�˾�~,4֍9���+�P� 7���s1D�o�{��.F� ��(����)��T���Q�3W6�gf��1�Z����/�ه��7	¨���Q�qs-��<��:0D�F*_>�ge��/!�2�V8xz���E'^����r�w��yi�'-�����x��U��ϻ��,V�Q]���cxZ7��љ{ƴ"O�%M��D"R�x�G�>!��F;�I�a��YR�$���ÌaAƗ���
&	�ŪM�O�!No-�|%�R�\�k��֧|n�#I���|�*�B��~64hA������ U� Ʒs���+^=0��~,�K���Ė�G�$w �1��/�竘_6�Y�L>s�g- �=Ɣ!a��|JW�O}�j�|��9H�	��y'&���8�>o���y�Sh�ȄA2q&4��%�����j����<��`G8�ǉ*�r�r��H��p�
���鍛�߃>2=��9B	x�,-@����/��o�U��A�� ��Y%�BA����8�yFI�� G�vq�Zd�I�jf �7w�k�Q�=�Q&"Qa$9F$��=ǟ��P��?<ZC�K����\�Ԫ�F��(A��c-���]��T��ݴ�2�L㇋$�6�2�UT$�d�pѢn�R}����F���K����ՆH�z�i�pZ��3/@:^KqPaK��,hՎ�����G�A,��D"�>`�|Q%P $��#��d
�f�a�$!A7������y߫�۹��槾sܹ�V$zJ"��H�> ��x2�DK^BN�]s�k��:�9g��\.wu�._9���ڌ�! HcE�`X$�� Ҝ��.�ߥπ|8���Iɑ�~��KA�af�����>c�q%9fYE@�J����s�3c=�2}]�3���3���kpp� �4��h���G(����8s����-��R' �䦔�1�6d<%�`�����8� �(B,��%��4Ꮛ>�����黝fc��r���I�=Md�� ��[nC�n���35a�Q����Y9��H�g+�[疰fs��L䜫NIG��InA'��mr����n#FfqX�%����AI�˸ɘUWbv�X9�ɥ��b���Z�C��PUHdW������4j�ӭͺ�,��^x�yM�yb��DxX��Ä( �1/��Z0�&��f��Iջڵ5Bܒo.̨%�lN�ЪW5.?+��Gp��'�c�����A�8L|���Z��8��o��շ��ݩݸ$�a��>qaE4O��>�g�-Z�"���9�]R��X�/�@>�F���@��6�E"BP�C��$͆F{3�LS�a��Nx���G-�`�Ò9��H��o��[�|`f���O�r��'>��*� � �N`�����Iy� E#*� q�4�$F9�.F�Q���z���W0�@��(��y�(��<S���5px����xf��� s5'&G�i-�A��s3q8;�lB��A��<T
>*BP?��s�O��bgw�|�����������{1��Ü�t�L0�����W�;���3}�D�"���H>\�Ғ�sm���oq��!�����E6d���4�	gs�sFi�|{��QW_��i��|9V��I��SY%���C����=�ϝk�}#c�"�ֈ���N��E󒮖�A�ͬy|��8���r�1����k�`v����xx@���$��̓p��^���S��߸��hl���7p]��I��h��&�3�>���貼��c^���F�]�n�e���zB���!v�!�`"0����Vuκ:��|ꭜ�Z��qC�N� �H���P�Q��MI�@�,OwbbU&%��n�3�"=1{�0}�@�V㾺k:���1�$��(�NfH<@�I����e�U}11?0Ͳ��jrO��Kp�=�����a�0_y��V0È<��XZ ��$�H*ӔQ�pj;�������<�A�m�H�A$�紃Ls��7\��[Ӊ���ԙ9R|A�Z��Q�-u'��u������"�&I�����8�g3nȷ���Q:5�A�8�,�� &$�b8`͝�_omtM��p�i9�8}~-���i��`�0Vmz]�I�(qψ��%�w4���&��{�8�4_%�?)����:�8� ���K�.7|'���\��e����aҺ���R�*GV�};����gC��M�K8�]�Wu=!F3c�Ů�N�Y��������Lt�+�m�Ad�e�;����EVlچ��H�[yH�ʼ-�E9ٻv-�z���O�%�K�B���"U {ΝgӔOe7m)CWWOj��F�xe��W�������w!Sp�A�@�[�Kj�Uǎh�$Z��R>�w�{1F(vh��ec��b�Z�nkŻt��R�G[��.Εӹ��B�d�[�i��%�v��=q��0���a�f+�F�u��K�5��{D�	T+TT�8��\��^%V���C}�������M#J�j��ҭm��O[]&�X��r�D�嫊�qy�;��O(�j�I�W�^;����޴c�RY^���P�$A7qT�Un�4����|�thɃj�R0L�Dn�"���Z�Q��>����������*י�w7g�Q:qi[ON�mfNۂ�d�0!�fҚsZ�]���\�0�sj�SJ��L�AdMItԾS��U�tB-�s�6�
�Q��sHQ]{em�L#{v*;*����[��|��צ�Y�,V�X��Y�V�\
-�����3�	�nJ�b���sc8�I2�ꬱ��������(ֆpG�gn=���x�u�<�w���\��om�m���$��nݶ�$�[��ݻm۷n�I.K��I$��^^Ir�I$�I$��m۽�nݻ/}�ݻv��w@���7wtn�����{�?��]�#��=��M��3 ����<}��h ��%��Y/d����p�B�A@6��K���o�s�3(Aӱ��o[����U����+���妋#^���j��Ru@�U��b��Dw���ZI��4%��=�����YS-9]����,����i�w�^�!���^��{�3�%#s��0���op��)���ʹI��B�̻xӜ͛���:��;)ޛ�
��6�{���{[JbШc;̊�i���	Ș�p=隨k��ɷwt�;�p{ՋWR�jK+,S�1��֎����[n�����c;+͝�Vf�)�.!�'-q6���N]�Y0��
�Q�缄��[N�����\�j��Ǹ�e��ʓdk��Zͻ��5GU=t�����w)#���qX��g>�k�:�]N��F��	�ג㺞��wr�D�K�m��S��������E�0Z�t�o���w��^�*n-����i[se
�y4qܝ!y���K�K�z֎Y��� ڨ�3Җs�5�U}٫�WoX��B&�^��J�N�q������0=��Q��v�ni�D�qu���l�mG�f��1���,��j��8=��U<b1�Х��wR�T�{�y��lT��]9�K��vF�P7Qm��^�J�!kHb낁=���\�d���Jp��೹��sMX��t�˺A� -�wQ�S��djR�}A�ViG8��E��"YD�B��Ć=�wq⦫U_3�wiҸ�8�`P�E���b���C��)y�4³�
���D-\V3�^a����;�u�3.
P�M-hK�b�i�ǣ'Ng:5I��+5|ő�3X��ݑV����{B�ZQ�f�u�P� ]����#C�`/P+�Pe+��$���d��:mc�<ےWJW;��/�����s�t�Q�Bub��L,݈�r�<��i�]����/���x�]"E�7���|&eJ�w�o�,�-�+���Y1�s�1�(���vKh7M�Wok7kŹ+��)�|zA�Ӱ�2��#[`��4�����MG��n+4�G8k�vi_�W��
)�c��50N�S��\��Ϊ�vs�F��N�N���1z�V˾9���v��Η�L+ʊf:��u���CzBN`޾e뾏-9G�\��m��F�oyNu�7��K2/-��r�ן<Zݮo�^��fb�+E�o6�͑�`,�Y���(�>}t��y�Y�ďBT��>[�H�7��
MI�|ptb�"jM
�(�$�q/z��q�xXCI���'A�!�/	�4,����w�vDG�aG�_|a�E�A,�iNR4�H"0��jq<�cV��Ҝ:鬒�D'�8�F�������Lh`��?�.B�aX|IZ��i�f ����o�/s:�A6�I�@��	,��K�M8a6�y���!�!Q�qZr��� �3�}�T�\+���iA��C�9��I.9�A�9h�(G��������g��Oj
ex��(�Ě�p̈́�K����F��D#;��8�d<Q�9�rsS�EK�ƃ��L��&I�AbNL�qK�`�XfNGQ��\h�ҝ�lV>��ȑ�cEfl���/����cC��Nw����`���4`@�1�w���I�o�Abn�Iov�}��U5׹�����0U��6v��)7j�F�"Zf��v޾�M�y��ELXh�h�- ��axY��H���qJ@7L�Q$Q��R�y�T]2FJh�cq�AOJAa���>�epےKI�ğ�,��#N����Ǻm��R@�*w,�K�NQ�c[���*�3'�Q8�7��&a�$Ih�s1W���ާ̋�����#�f��Ϥa�p�c���S	�_*��h� �| ���|A$A\��7���T�Oa^N��$��qG�`�h�G��z}vW����.B�qZI�"�9Em$����;�;o�pǐ}�ɓp$�G(A/��Qv�0xEd.�Q�,B�aZr��$��=��wg��D.S�Q<9�x�Iq����r�����E���X��5����r�	r��)6G(���Qvj�X�� �����Ӛ�f1[��+W�����󸏩�����)�ac�F�Gǋ ��(���ß. ��=GR���9P:��.ݤ+fUeUb�{����O{B��{:�2����R�<�)i=
+>t�ORb!-�ȇ�-�Q-�Y�H�����8�Ay��hB�iQ�<	'Ա�H |O����V��k̶�������Nz����=DIh�A��rHFs�U%���*�g��!�OAh@��(�c�Q\�J�����le�qn}D@�bNL��-�Ꮝ�a{ۅ�ߙ�A��8��,��(�x��K3���������0�ɤ��kpp�=��gȦf��8�� �����H~JD�#Y���-���+�s��I�ne���gI��0�����7����H,� �E#�r�'&����l.7�VLDT�ǚ�>At�Q��0r�d紸8Nm���'|f�|%d�Q�*ӔQ���[��'#����*�m����K�������&�+˚��R8����V*!���qQ�=���4gF:���.�L`B�1��<�Ȃo��x����O���̹hY�n^bxgp���V���5f&�:ެf�5Z�4N�UQ���9z^�����)z��<E#G��>+g�Dqً{��>$�IxĽk�
w�DCR`�ãZ)K��:$C:� �ӂMNL&hT�'��h,q�	L$ӎļBCZ��ȫ��F��6�r���+I~�xH�8PB\�i%ۄ!a�Qc��Q}�>�C� ��Q�Y#��A�$�I��^�5/��K��� ��D$��I�U�8bJ.��Mw\�ߛ��A�&�Q�1� E92A�p6=g|��}����Ώ q�0�Y�QC�iNp�|z��&1��$��"+Rrdp��[Ih8=�\z}G��� 7J$���>���F�!(E��Ĝ�k}�}���긾f��Ԝ�� Ʒs�4�Nf_з��"�~f�(AC�Y%���%"rF�JM�OWGġ�Ҝ�g<�o�q�"�,H������k	�dy\fl�ʹ�%�O���U.#6�LMI�<�7m��%�w���1�O��iEwt�nw���������M�+�W][����W�Kq�5w	��;r[�OhX��@8M,��h�K��˻��]�s/F�WR=��3iU�G�x�3��xYUL�m'd���7�ќ,2*�"��0�R�Q@K���^F�SG%I#E�F�h7��Fek�k�����M��0�6��)J �I��KG�7oq����ZK@�<qE�<`��ϴ�)��|*W]�n,KOQ�*ӔQ��In�������B���<����(s	p~É.� �$�H8o����z���(��ӟ6$r�3Ě�ac�K���QV�}�A�AŹ��I	Ϥ���:�4��H+���o���%E�I�@�,rd6��-���{�����cDt�⏄Y�YEA�&�4�u�ex�"3rdp���K@�x�N���V;���,��Q�HJ�y�����.�����q��;�w�%G<�5��v���5ϙ2��ދ�	Q�¨�@�X�0M�JԹ�#8P��`�0���Q��]�0@{Zn�7��.$=S�י��h�\y-v�L9�y��k �l��	�%�;�Û/3�{�ҥ���0‎�����~�AP�-�Z)��-�)2�ʦ�d>`@e�"T�-4���Z�n�z����NY?k[���l�A�AB	��[�>5���wSs6�K$��ĤNA�i4���m��7�տK�{b��
�(�"�(�Y���8k4����^Ǘ�4�~��(��I�=Md�� �f:nv���9 �4r�d���)�������a��K��#�NaF[I%�D�yY��E���0o���m�A�q�i�(�/�'��_}���w����Ü�A�In9'ŎA.9�i�~a����=GF/7ȩI	ʓ>V����8�ѣ7��DE�"�0�$�h��}xd� @ ��0�C�#1H^)C�S��¡�\���`z,n^�"7�z�3�gSnY�ɋE��]�$n>w�,uR�$�4��(�
>,���s�ӤQ'݅	Z�C^�S�ݖo.�{�-]î�����ܥ,�����|RVE�0RڈI�s��B��⦄CyA{Ђ�>&��i��C�>�5@�.��'ۮ��}�����8Pa�anYEA�&z���a��/s�5R�`�I��p�����8g�i�`�0��\-����I�Q��%ع�����&��v�s0���T�G÷�5ʓ�,�(A#��K� ��1���^�"8.$#��4,8�G9�U�^�U:_ �����8�	g���PF�H�s��r��z�_6�q��2��-A��Q�F��G,��T���p�ܐ��!� K	4�DU�8c�N������:�{	���.	>9Y��K��I�5b^�3a>p��H$����9E�@Ⱦ���:<��/.Q��(QS�v�N#nz�����ړ�@�{������D��;���؜�!���-j\��u{�1}Z�����_]��j���1��Z�����v��㪅����<�^a�W$�R�/j��{˝���H�x�Hu�H �S]��&�T�(��]+m�Hx���H�I>�>T�;wfIe
S���.��A,XA����Lr��ͅ�t����̛�lԐ��A�*��Z%x�\��0�OO�)`P���pZ,��h���ok}��c�1�$��,�	�	=D@�bNL��dZ����{��Og�O�8_�$��0r�*s1R@�l�}�o(>@�*w4��NQ�A�np��%��"-�\�,��0��?$�R ��73v��;�Ǚ��!||9�4�������gI��s?�����	��Y��D)�D�(
 �G�Qp�t[7Ҝ:��Ih"��a��)u�:w�����]X�uŭ�j���z��6L����
��˸a���q�;�s��{8�#ևP�2&��o��+�aQ���S���oo'!�V��7���qO�m�H\u{��n���vj:jU��Yܗ.s$��ҊP���շ�s+eռ�%3�D�z
*=R��>UO y��Z��'�"�9Ed�N���=����fo �=�>D|9D�?�i%ۜ��E�rO��Z�`$�
�0È*ӔQ�H�v�q��\in� 9�9�9���A�Z"Bs$�r
�{���=fg�Z@ei%�Q�>rHFp1��f�s`x��hИ;�Ah@��&�h�1�(�f}�-PC��1Y�	��:���Ԝ�>�-��f�N7��z��#F�@uIe�Y��(�x���<|�����f-�w>$��&��}�5�8c��5
�׏L,a���4�
H�Ih�AHDP噫�q5�آ�����Q������1��:>����Fv�r2����k�)�#��*/f���R��}٘��.yH!�c0 �a�%�缒��@�a�t�Qm��E7m4��$$M�M4�=��7z���~*��p6�̪[3y0ę����G���u�T���s�}�A�m�k��x�B's���#��3��9��ZA��M(B,Æϐ�u�yw��_B,(D��L�exD�pݣ�o|K}�[ϙ�G>AL�qc��*R����j����<��c7��`�x��U�(�,�Ip��ݙ��7�
߁�� ��"4r�px�K� B��3<gu��fb|7�A��(��Y#��A�9�$Ꮞ$^Q�[A��>q��1�DBHNg�<"ih�瑻����dI��Ad�9$�&C`��Q�s���<� �i�,h#�e9��]�������wt��q�n�<�<�����ف�M��덶�o�����3��6Φ��-�c�Ń3����jٛ��l6����������3~,�6�m����<��ف�o�l1�����Ǜ6ف�������>�m��x�'�{��������m��b�F)�)��51L)�6S
��LQ�1kF-�ń&&���A6��LY�!����&, �1l�i�i����M�b�-1�Ę��PQ��Q��
0)�bALP�L(�P�Fb���0�l���1M�1LI�1i����LD��1l���[i�� �����b�a�3LX�4���Aa1a12b&�&-�&L[LY�Zbъ��($e��-1L$Ʀ�LPSbM��1#aALI�1�
1 ���(Č���і�&�i�h&� �1��śM�&#&!�,dų&�&&2b�i����Ŧ-1h&��13&#b�h&2b�Y���)���Q��1&��1LI���$�1&-��-1M1db��LPH� �6e1LZ4��b&((S
�L��+
d�F�2����,͓,�3!bm2i�&Z�#(H��	&ViY��e2�$�L��mbؙc&cB3&[m2ke�)�ȶ(Ze2��$j٩��e
�2��Q��dX��$�L���Й126��!��fm�8�m��m�Y�F�d�e�dX��#L�!l�&&M�&&XB�L�&X���ɖl�#m�C6!,�	�f&[6B�,C&Y�5�&[2��,�d4��F�-�d�ɲi�F�X�L�B�e���,B�e�-�!bB�Йd�L��i�2i�B�&F�	��bdk�d�,�#&L,F�#d &L�2Ͳ�1�#2e�ɖm2ƙb�m2�2�L�e��L��L�,�$șm	�Mb����6��!	�,�Й2i��	�-�m2ؙ6�m��ɓ&F�F�l�6�fL��12l�cL�hLɐ�e�,�&[B,m�#m���[X2e�&�e��c-�4ɲe�2�2i�[�ɖ�	�ɬ[&Bd!	�X��d&L��!2��bdɖ���e�ZemF�)�L�Xjش�	2�,S(S$�F���&Mm4�2ɔ�mL�S(S+6�VĄ�-2X�2L���F[L��#L��4�m�6���&F�&�i��ň�L�ѡ�be���!�-2 ��e�KkFQ��H��L�[e1[6�)�d��)��6�Sd�jd�B2d�ɍ���2i�2d�Ћ�$�L�$�ئ(�S	1#mLHĘ�F$�1 ����-LZ2L)��LS���&"b�PSaFh��lZai�ALZ	�"bASd�Abd�dŶLY��m1fɋL@A34���`��l��b	�A6&,ɋ6�̘���ɠ�b&"���!1h$�LQ���m4��b�D�&&�A4Ŵ���&��&,�ɋi� ��-�,LBb�6���bd��bi��b4�&,Abb1bb�&-LZ	�,����,LM1 �b��LD���FX����LI��[AŶ��1�ųLY�4�1f����[LF��A	�&?��߯�6�0><?������l����|?���_��l������ف��l��o��m���v�6�0?���t����>;{t����l��O��f��q�/��l��m��������x����:6�0:x���?������m�`3�-�l�����?�b��L���� ^� � ���@�  nO����>��O�fiYm��*d{c�;7�Z�<USlVCi�ci�4ՁY�2)��(�Q6����צ�+6TQ��o��        $L�1�Z�5V�`�!�i�m��̵55��֭�����Z�i���j��-3V�ڔ�&��lU46�cM2�i�f�Z1�Q���-�jRֲ�&���[$#%m��6�f�Y�5�ͪ�U��Y-ٲ��� ��ka1}���Z�F2�4�akU�|��y�y�]�ۺ��q����[���v�YѠn�Y����� �n�ε��� �&C2�h3[�;�жmm�e%TE���JR��)g��=IT�)R�TwJT�T�[�[�J@ �3�T�7<ۀt�;� 6Nۀ 1n��5��� ��T�نK����D+[���G�S��kU�J���\�gG�p�V�vnh ������@�`�v�Y��t��SZRO �S�Zm3Ph�V���S�f8 ��� ��s� ���5Ӏ ��� � �0 \�\ �I)���o�K�4�KH��(��S� �T� 8f ݎ 9�&!� �q�R��w��� ��8 �0 wAE�M������Y-F�[m��Z�@�e� �� �׽�� �gp m�� .� 3��� 6sp �m6o��u��6������R�m� C���� 3�� 4X 7v����` F��� ��0 7 �al����7u)�جʒ�j�6� պp�ʌ 	�C��#�� �sc� ���� NA� =�gH \�p ;��(L�ݍҊ�&�Z(i�B�j�� ]� h` w]�� �:� s��\�7 ��� n� ��}� w{5��@k[|�=�z�	6&m���ER��w�z\8 �p wp� �p *�� �f����\� ����p                  �T�JR��@�S��RT�h&�	U1��H�UJdр i�S�%R�   ST��OD�I�F�	MM�*Sj���}���SJ��?���q�8DD� ��!A��ޝ?��f��Ѷٰ9��a��m�`3m��?�fٰ?��́հm��[6�`�c�?���_����R+����������)�^��M�\F�88�VIX�ոxnb9g���!{v�Q:�d�f+��a��-_u�f]kG �K"᧩�>��j[d���a�B�M[�[���Z�(v���q4l�q�h��Wi���UK&m	I!k�	����w�<v���і�C8��*�]
�x�,�N:B��n�$�Q�e�0���@��6z�r��N+��?21�A����$�a��!Vk^X���(����l�8Q��j���$��餼=dx�]o��.&$���Q7�a��aknV�Ba�{PnK���Tr��+m���(m:��:��f����A��]Szn�eS,���9�X��z�0���ECSEy���hӨ���]��^Y�.�A�l�^5��@s ��1��,��e��i������yZ����[$絙�D�ܤ��
���ؚl'H%h�%��	��n(���e����<0���0���$��ŔYʸ�eZ�A�r8��Ug7����y�����0��+W,U�Xʓ^�[�mHoI�Mݫ���Ě<bXVe^75ηEz�]^�N�̭�5:P;9K*�e"�(�[�CM�K�����2�Ec�����:ͦ&T���p�ow.�P:t��M��EJ��� Σ�+�go�[F2+
^]qz����<����y�^X�u�*7VՑ�Y�Yb`�sFcF)[1�ovn�V�Z��]S��n�뤳eR�Wy*`�c!A���ZS*��}cxҳ�3�� �-���n����3U�k�V������S��)
�,$a�B[���_��cMnnn�����)XU��%t����7E��UQ�Suq?*��$:a�@� x^���oP~e�U�̉�a�[U�vn��{xe�[�7h�b4����Wђ�n�t�%��6w"[W5Z��Ȼn�:�zUdK�w�)�K�J5��Rbӎޝ�
Ï[&�a޳֐Nأ�ֱU��g3���%��b˴"U1�/1�yI]Ih���E֭�V^?;�VU=~j�6g`2�E�>~ڸ;,bg�d�Y�)���ÜX[<!Q4.��]˺hҼ	2nҒ޽&V�r�׵cV��>���[X���N���s��+.�=AM#Umb)���͠sP1z�Ԟ8�L�N�\�+���=\,��Ey�C����:vY�-�2ࢋ�K+�$�h(sP�d%�T�4�="&̕��_�^f��dn˫�w���*����z�lRN��n���Φu3ɜ���L�3���#�%��}z�B��O�N,���8�y�<���%����v6Beq�f��2�u	Nдj���XV3lS��hVk��x�!
�Ͳ�n}�b��gD-���h]����ۦ�,r�Lr��K:;뾣��}��w#��	\��Z�z��i���V'��r����=�l�s�bhټeb���yjTM�Ecyҕǎs7b^�e�u��*�v��̌�5����X�ωr)Ǣ�n&�����t���r>]����+N��[8��'�ۚI�o\�2�v�g2��~���څڜD�Xv�*u�iG�#��dxi��h�2��s�k�TAGl>�����7i�N+ 9E;��"�w��<	g-���Φu3��s�:���˝�|1_	�^���o��U�$�]��4Wb��7��ō�4X3" Ԭ8c���!j	���z�*�;��X`%��T[���W�7�ġ�Lš�C��x<4�m
�6j�7���VSO`�U��zaX6����g�MHJ�ѻשr7MU[b��W�bW��jru����"�{m�S�`�3��%�)�����C	yZ�|���P�Х��%��k)���n�咒����1G�Ȟ`x�wnɑX0��ll�%Dv^��xB<,��9Ő�]QJ�����u���suAR�8���hF� ��Ò�x޴��T�:w�_m���Q��EG<=�23�K4ˣjC��FUR�hYR���N�u6�$v���-Zn�q�S���LK��^�H+u�S8�gt��a��;bj�r�+�]QھM��:^�K[�ٲ�ڴ�q�k�Q����Cr�0�ݎ^��t�u1(��FhO��Ḱ�+Q�Ǫ9tO���i�����D�+�Ԁ<�hN��Ƶ]�ھ���\c��Vdwfot�p�[��v�AL��o[5��< �"�8pÆ�$�h�'O0޻�P����đe:p��͛#$�Fh�*MP���0�Q�G�ae�C0��{����%��u���:�(��-T^�KU6��ˡ#�$���e�7�o{f��GfZ��r�]k�͖���G����;7egsl�z��JW��/q��Y[��M���!";�퓺J�ڮm��(����m�tgI{.�}+���������0.���v�K��|���+:�	���ԖV����gf�8Id�(ٺ!Xi�&�*ĽnI��#����Yʬ�oq�#zw["�����#��i���7]N��|P��fbu0���fɭ%+�:v�rW;���Gt;|W����/b���f��%�ާ,`�}�Fk\�ۢ��\;���zbOE87*��B�����l'�S=�
��9�ܗΪ���-�n3��nVd�Ai��S[:r)ӫ�0�BUv��#f"�4p���cyC7�Q�� �I�A}�YX����}]KM x�oQ��O�37TVX�WA#eEmm<�b�,4Y�m�o]uq�R�mO�Bm)��H��K�4�k�g�h��:�Wk^G]�g�L�a'B�Y���_G�WU�#�i��+���st:L\ˣ9�YdP�4G�u]'Z6���3�7�)Ǔ�
H�Y��C9�]��Rom�6�V���3u�/�Z���9y��u�ڜ��c9� �7*�9L@�Q�_Jٕw��]PBXpe�iG�ݬuy������v���g^�K�7g�`Q�D��S����vv(QN��+睕Bo�S�L���b��dK�:��̃u�p����x�=��YP*ذVF��
��T�JKM���F<Y������ʫJ�Oa���Y(G�e�H+uJސf��5k���o�ˠ��zcx��:l����[��׌VZ�O��g�<Y�)ѽ��3*Y�\��֟(�'����.�a�ܱ��]/R��$6�Ј�n���f�Q4uF���r���U쳩�jn�UV�W�ݭ�H����m�vS���9�N]t�����{�kK�r�+v��bP�g#m��5BlSr�6�SN�,��h�LmRab{K.�iɤYA�rn���Ӂ���+E�)%1ÕԳp ! x75v�(L�Mz]����]d��B3ם���;9w���c�eT����<f�n�6.���&������ՏB�gȒ�cyV)c��r�LeNS�'[z�� ��{wj��_+�W�O&rp�s�d��r�2��{�͉�.֢��v�W
�Oy�6S�[����Ĺ�k�j�DGr�e1�	}4J�A���st0��p���y���'���@�D xQ �!�F4q.�'�a]���!���jU~q;r���+ܫ�F"$�}��7�ھ}��a�y,�	�n�S��5Aj��L�T��4�Z���(�\�]kj$�FȆh�K<p���p�"�:a�5&�!�ј�}�;���W�CU�-�EE��&9Ztm\d*�j��1���LZڨf؃t�q5pV�]���.��p]�P5�(���Fb������D�]yZM��i0n�q�|<�<8��O��J���$$�)ʂ���|
.�
�w�VQET�m��l�JE*�ʎ�Tnf]��W��!�<>�y�g���>�Q������a�-�-H�[Y=e8e���ѮX��ǰR�#�N�Q-*�m�]��L$�N�/��U��={���t텻���4�c��KE�@+Ut�b[z����J�C@�:+��^x[�h��`��x���)�&Q��mRѷ�i�i�Z��z��%��0b@�{��Ƭ�I���ګ7NZV�J1jڕwLH{UCJ�-kv��[��Zm$Aɐ�*����=B6m4�
s��o"�e�q�A�Εd���2`��E[Y�"2���{-�J7P�3���@�� xB� x#	7�{��V����X��_��;��n����ܵ�@p�]+qT�z�u��`��tMa�)F���W���e�Ro6&�b���Ϟ|����o��c<����3�g�ϱ�F|���3����l�g�Σ(��<��b xY���� :��ɦqv2�����8���iF�x��=ڭ������ˤ��%ַ)�{�n�&E�!��a��*�e�fSZ�l3f����E�34n㚻[���hZ@�J���j��a��gf��޴�Ub�IK��k����6��S��o���GJf(/�[�R�vB��$u�a=���t�eQ՝������x�f$�C���6�J��/0F��U{�c�<��#B=�����P,g�L.E	��B���+����_&CU��\�H�������|�R�S�#�(��Ma�@�p���n\�u��2r5{�톶�+��y�(j�Ò�Od�>�w���o#yh�1#L��i�	\Sw6�qK�b�[����o���c+y����0HW�7���U�u��9��km3XRj��+l��oV���L�v��S�
5~|�����ƅ��ˬ���;��n����`nk�CF���!�ir}:�S�X�j�*���<��=�n�D^�W'"�	M��uRi��auϹ��;���z�o�VH&�h�C2�����]��"2D�r��v�р�Z�&�$���
s�!��U��qJm�̊�<Qʯ !ҋ�g�\Y��+I\u�v��q��rh�T9�P�Nk*��4�B�Z��8�=w�g}�q�{�ԷU�x�9HMŌ]���%n�J�cF�����oۅȋ	zQ��T��8�-��k�j���o)Պ�12e�xK�j�Gf`K]*�a׬�V(��v�.��n�a�VQ�ea$�t�/�S��Dv]i��jǍel}�I&�n�NAݎ[U��,�v���(�T#�i��(��pCf.&c�3��D<����@àb�@�� ��wm,éT���9��GM��U[�v�S���d���A�m�a�xo4I{�M٪�u��4������	PL��0拱y����x'Op�),��}��Zo��Eڝ���A]�+�N�khPu��5Q$!y3������+ ��i���Iǯ4�[m���\Ƅ�U|b��-��k��!�q�U��`�\�yv�5�����p��7��D�0�F�� �6�ƦR��;�[A^1��`:w�R�Ƥ��7Q�vj�.��}�f����y:<=f���#ۭai����݈a��-�C���c;���So�0�+a�n[�Oo��;|1o�9���د��:^m3���IW%��f�8;{�g}���A�UY}���q	q�k�c��u6��3�M{�)G)�v��*�<�.��^_�w0t�ۼ2�N<��˨�N��<(�o��6n����d�ݼ���8�v�{y�'gGGp�·��Je�ws�t��,������ߴr�����6���ص�'}dd4/����=#����-�Q����٘1;�u��L�g����'E�u�4��x�o�T*�$��J�q�9[�e�l�9E����Z��g_ ��h{�m��*Fd��}�I7����i|Vm�n�sCNY��!�"����E�� �˄�5v�Z�E(��sC��SX�v����d����0���m�j�ˬ60j�Z=s\�����X��&�f\B��)�"W.�IA΄	44���
P˘��/X���hK�۫�;8rܟ�J�2�^+��,-y�Ir�c�t������O:���+a�����k���i����T���v�
���زgM��l�q���b�Y�!��;���J�0ڎvd�.�i�E0�]| ,�IP#2pم�:`�n������b�_[(�]�$�����]��v�+�퓧Z��$4�JIm�7o7��w[wiem�K39"R\�K339 ����;����x���	.�^I! �Y��Y I$�^ܽ�����I$�@� � ��I$����~�0��I-�n��I$�I$�I.�^I$�I$�I$�H�33:��<����}�:��@      }��    �����s�7xff`>ηwC��{�gl  ��;;���}����s33����3<�nffs3ww�n۠<t��������vv�� �: ��u���}�>�κ�  ��h   y��}�  �30 ���    \��ww@  >��   ��� �ߴ}��`      u���  y�����ۙ����nffs30��g����7B ff`733����m�Yd�Kz�,�I$�,��$�[�Ye�I-�,��m���%� �;�g`:{�f3�w^�fc�wtfffs����}�I$����m��$�\�,��$��Yd�Kr�,�I%�{˗.Y$��Yd�Kr�,�I%�Ye�I/���n�It��I$��I$��I$��u$�Iv�rI$�^.�$�O�$�__O����$��e�Y$��,��$�[�Ye�I-�,��$�wm��{{m�I$�,��$�[��r��$�e�Yd�Kr�,�I%�e�Y-��<]�������o.\�d�Kww�v���3�{�{}e��˗�]�ܒI.���I'�I%��I$�̲�,�I}�Ye�I-�,��-���ff83�<���������I$�I$�I%̲�,�Is,��$�.[�m�I%��I$��.�It��I$��I$��Ye�I$�]I$�]�ܒI{u��m�I%�e�Y$�ܲ�,�InYe�I$�,��ws~̲�/;�{���s\�m��$��Ye�I$�I$�I$�I$�I$�I$�m��x���s30�������o/.\�$�I$�I$�I$��m��$�I$�I$�I$�I$�I$�I$�巶�$�I$�I$�I$�K���wu$�I$�I$�I$�I$�I$�I$�I%��}̾����I$�I$�I$�I$�I$��.�I$�I$�[m��$�I$�I$�I$�I$�I$�I$�I$�I$�K�����od�I$�I$�I$�I$�I$�I$�I$�I$�I$������$�I%�e�Y$�Io�����G���)�nbIC������ĒS33*�$�I����T�y�$�$�A/$�y���q��� ������I$�I ��I$�I$�I$�I$�I,��m�I$�I$�I$�I$�6꫻��)$�I#mȤSws32'�@ooo���Y`��|d�$�j�H���6�}��#vX���o���A�AI'��+E.����j���7�Y�8K9��i���.2{9���]@��(۠�#�+��'VЭ��𺈗sy�.�'Qm*�y��^��[9c�gͫUW�Qm�u�l�^R$$�� R�'US��5��D��2���ƈb��p(�S�wڮ�,�{ؖ�]�
[;R�:�ۂմ7�+X�����az6��.v@���SMpו+���6�7��-۱ni���zYUºa۫������z��k�Κ6�����D�������UB��-�-�
t�ᤓ2�1�f��ӷ���D�y��
ܚ�w;���w�Ҁ�۔��[5�l-ŷ@�т��w[$�鏞gp�p�dP4������c^'g��J}�!�K6�����-�f�Syu���˕[�������mF��>�
���ȅd|�ˁ�v\�Z�b���>���&f�&Ի6]�9D�lu㩦f��}��]g�
؇	����^1lmQNem�����T��J[R�j�ݗx���hr��� �Z�T�Ò�>�J<�*×��*��O�Q䳊�mt���!�uj�I5��^������v����&ܛ�:ݹ�vK���Y��Uq�Ӂ�fqYuy}kz.��i�%��\#އc�uGs�^�y�܃8L��4�˨���67	9M�n�QV�˫y��wR��lnw+��.Q��Dt�tһp��e��ۥ�j�'˸�{L�q�n�%ة9J�KD2�(�SZN!>y&Ͼ��>�b5������=,�${��v�L�z����xrO���4+����F]�1�=��N�z�U��'7���gsp��-�I�"�ڡ\�	���v���tMC��S�أG7�o�����&��a��c֪J�T�eRN����9-.c��_;���־�%#�X�K
�����m�ɠ�J�L�Zs�[{,'9�Ue17B��\��JP�4 H�+��k�.��BiS�B���ϰ��*&wht.7�+&��c�o!G�[�4�F�<��u��a5���A�Z��ζ,�|����m\��.S�J.�\�T�(ͫ��*p�ؗ=��k��:�Դ�TC�&rTUNBBƫ+6r]GJy\�]��Ttt;�ލ4U͒��Fk�ׅ͔����/��]1��Q"�n����p�:%kSz"R5�����ӈERt��V4�%���kK��g�m�VL��0<WG9����y�*�f�h��X�m]���U�ײ�B��4gG��.v������eVo�b�dl��Q�����7}�U�{pur�󖅜�"(�Ö<�{�$��;���7vD2�WM��aG5���5��!L3-��̓�י���M�o��k�t0u�㎷�LVf�.���g&73�
�I���$X�@���������4�ۼ�ɪ
F���[.�cR��'��[>�R��	��[��8lʚU7Z\�n)̳
�+J� j��K�mӠ�^K�)�2�@Ws�t���b-���W(Ê���$�gG[��K��r�����t`q����ʝʋǽW�6��n���vs1S�*��<dK�2A~.�M��]�������ky��F����7��xӴi�QT6ƣ�Ӝ�w!����7Ϟ^�Q���B��v���S���e�)���VJ�����L�G>�\[Ol�R�-�v{(��M�5�����%�Vz_4�1��V�ֻ���L��:�*���0�����in�J7�h>Vu�7��V�R�0�Wl��:�*�&+2Bk[�QÌu�RLG8�Z�0ҕ��U�:�xT�I$2@�e�#q7	�e:N�"�q����V���{�����[y�A7����% ���4�ᒝ����\�`V�C�k&�\��J����sE�zwp�;�Z�EYr�-e�.�'A��U溾��6��Y���em���tͳ��g9�9�rD�vk�s���d�u[n.駧Q�.*ꫩJf,��s�M����*���9椨w^�l��Ȼ��Ŏ�䒔��;���/�X��l�>4>�O�Kii���k�T��q0�N��*=�;�Yӥt�j���d��Wc,��H���\����7j���J�*%�$w�U{q𩝛ףyl�\{5U]GŲ��UUf��Cw�/qB�����4��6���v\�RBnJ�\�[p��5�v�؜����dn[D̙���J�ꆫ��7wm����m�/����(umK+tE�eXMr�ZC�`���&-_
��S,-o5�kyȲ�4+���BF�p,og"�C/V���q'���p�N��a^\��5JG����&�˭͎UM�7HX��#��%Vsު���w7��A�Z�f5Dt����-�ѽ&Ɏ�ATL�}��j�3��K˻�� �/���iXʮj)��YOcUY�\0m��J�,��&^��&K�IhأU׊���2�zsf�mԑ�ȩ���Y��jzz�[".v
Jw���j��o�=w���B�;%wS%���ʻ�w��>	UZ���-�x{��-�������b
N�\�盜��&ꧼZ�E�L?�����}�m�|r�[�d����$���ݛ�4�ڇ��پ�QU�������O5�V�2�8>:��wY�3\��{�j�����&�ޠ�y�'f��)�>eN�`Ǽ�����nJ�&U���{c�z�l�����<o��|��v
x�;'d�/Rc�M]Q¹�y1�e�i��cG��;y]C�WU����%�H�����.Mm��q'�|��[��}�z��鋲��P����g1��f��8R�%��6�>�5���ZA>ۘU���M����,%���"���j���d��!噗eWG}ʅ��7cdV�Ii��Y�^C���J�^�5��k�ևY�v苮�T�[$��36���R{f�6�ƴ�\N5�m.�y����$i�/k�
��$͹q�2��X2��3B��sA2�=��l�$=�洫1�#/�	��;�IAִ[o;���v�:垻�L8r\LE��j�op����ǣ����f=ؐG,sXmC�r��{FAɛ�U:� �w�q��#K�7�ӆ���Ns%Ue_ɤ�������U�p�M�>�����E�e=�UqBf�wW��R�}ݨc�ϲ�H����,\�0SkF�<9�v�xm�9ʃ��o��TI��Pwe���I}ދ����\��Y}�Ō�[}R�`x�l�]o[�*��XN��Ct,��f��98�����*u(/�cPf܏7F�B�i���=r�UEO\|XzwWqأˉb��w����.�c�M�}{1�w�r{��v)�utI��R'�5P��Q�yЈiWp�zi>�۾%"�j:ͽ�wy�Zv=�7#"⛜��S�1.�B���w�gܹ�J�ned�׫8���8���u�V31^Ȯ�H�U�T���V�ɫz���Z�хI&�K;+n�[SE)	�vA+8WV��VV���$C:SƙH�ۡ�f:[����s���#�V������U���o��D�`B1���Z���kj��o�T��NE��(�'S�%��j��S�(D*�F�P,wX�O��xˬx7��N[��hA�4�+�ޥŬ�5��)$wsX8d�[���tJ�����u�Bc��*�8��v��}��Ø7��d+QΣ	m��l��{�Νum��o؜�+�uz�^n1���Y���Qy�����j�Zz�oBz�]>R�j��fI���$kE��k1LU7��yE\}�cՖ��7����7�"λ�׆�[9D��$i={�%uo�Ns�Re��M���4��L�3��Y�i�5 ^ob�5Y ��]UD��U(�ٸ�"�x/P�\�+t��Z���V�U�3(��5wq����;:�\�u[1,z:���:&��u5��ɸRPBeh����[�q���u{��]�<�(Nn�c�.bR��ߜb=�T�|WWW:�=$8�l�Wu���i�l�����w����b'����m��٩�����)�j>9��wv\��*mtФ{�d���٪e.�t�r5z��olj8ﴮ�����[�0�,�)���s���vU���v���l���Q\I������* 4�)�j��ӯ�@����N�ͭ���c;/��p�p܆�Lh�˳�J�K�]��b;Z�å�ݽ���u��(�m��Ɗa'�����x����2�ԫҾR�.�Ji���W������3*���5�Ī^�C���b\�,�U)���R�
�-�1��d�H\�2��2�,���(Hu����T�9�z�SƇ(S9.��LX�-(�]m���K׏>W�D)��IF�[��r��+��JmB��`d��i����
JQ��޶�����u{�h�j�w�BUZ.�[Ւ�j�r"�b���z�W,N�r��Ю�`}�nU�qQ�e{��ymJ\���B�]��Z��ʛ4�5.�I:#,$��|N��,�8���K��ⷤq��ٽ��:F��Y��N�xS�q�Q�%�!����֭��T}�9�ٶ��3oEy�b���%|�=�h�Q�s/ƕZ���#��_ޥ˴fS]�BR��RʱM��ZF�XX�سlC����p��uR�U� =.���r�����Lr�jYؕs8���3
�/$�;��m�0�+6�])5r��>��6ի㇜tw37j��]�ʮޝ�O��ť@g�6�*��cR��ʹ(*�8�ZSy�.8죇v�Ɏ��+���c����nv�:<xU&�g\˻���9�*����=s\��L���V9�][���5��6�{��Y��	7�Y�i�8�e)��pھ��R���Sf��dF)N���1���6�5��N˙Wz%t�+C�����#�=V�R]2�n��v�2��z�d�����h����!Ԕ(-���׻x�_=[��/��}��/6��/b�'Dz����ɤ����Z���9����]�7��2R4���Y]�B���h�mh=i,ۊ��x2��}�&S�10�N*;����jr�q�6�é˹;"��5ҕ�]pq�wXuao�l�>����ڈQ����[>z=�Z�g�H9nSp$�c���Aa'���hX���c2M�j��v��mq�2Hr�_m�w�B��V�8�W�N��Wc�v����u�����ѿb5�ٹa��tWwt�pͭW&���urnc[��8��>e=z���O;޼�Cn>«��]̐�HU>���n1�U�wU�C	33���ԝ�ҲȢ�!RJ�ћ�W6YH�h<��1`��ϽQ��I�ڳYۭݷ*�j3VT�GP�Gz���q����]��EgS�ؑ}M����]�v[{����}Q��!NfjH�M䙗6�J����/Y�*�����������o�m�ޤ։4�����D�<�ws��h�����
�/03mtd������P����-�?`{ަ��>�CuZ�wO����,�,�,o]��[C��&�ie�/=����3 �L�3 �'r�K����Yc<0ik�a=y����=��D#���b5����lU7Y�E]m1�{D٬B�q�@�m�ͼ�-�\5��/���W�:���<�h�������U��X`���\)���-U}\���:1��6��0�7��T��%j���13q��Z˪{\Sc.Q�TU��hz���x'Vr��N�jB�E����ЊH?:<U�m0�Ԋv{�9Q;-ؾVM�:}5�0@�}��zM�g쏹˾�W.�x�g�	�!��8�o.W*U^�n��צ9���S��3Bь�7v��|�)6���Z1Q�
���R�x{qu�4������,2`�I�D��Uvٚ,[�����!t���y��([A6l���U$��b�7�u���;w����D��#���`mS�o]�R���QJ(�ֻ	MX�h�ES���ƺ5.΍ �Y0[4�q��oV��U� �n�{�sXo�qE��ܳN�ۥh�hgw]����#Z(���o>�nc��b�����g���qL���7Gj����\�R�Ə�n�v6��k���#-�Z�0V<ި^J���nl�@x��1ۢ,�c��p�����Y�i�5;�v��f�ҘU�.��&���/Q�Z��v��0V�>����{��Z���t�X����+rv&,�����y�4:����Z��A��
���GK�Ǔ�n��'1T�H�J�o�m��Ok�j�e��^��CYs�A�<l�;Z�,>���C%�u�FPh:3j����X��7��M�ܦ��h�����\��)yk�j�j|B{n�ꮷ1S��ۓ�-�ӕ�dk�\E���ެԋ]j�]KxQy���U�u�/vHm뗀�αr��� ��4i��P���K�)���]�'.�t.��p̏�E��2Pul��lyt����='Ko�ޢ��NB�,��gN��v�vK�y]y��z����Ǎ�(���m¯o���KU����^�k�܁J�};)T�}��;<����W�_H5I��RC:�)Y�m����>2���W�ö.35S��J���8���ɉi����ʾ��7^\���%��J�.�ݧbX|&��N������W�R�'�&����]B)��͝u�����u�;�q�
nrm�N>YN�y[fF����L���j��ڮy�mn������QU̦��]�.і"k#+LZ:��,Ezm�\Sۻ���G����+V�\�Ԑ�P�
:�IknqBC���!D��&�t}��R�Q	]dI�uv�Z�+\���O�B�f$��+]��[sT�m�HIjߧd�Y��[�6�2��F5j]��]�:��q�ܔ�Tl�ʻ�^�J�8�:=���-�:=��D�w5�9i�-�y�$��%�բ�R���wz�vCB�4%Ї�)
��L�MN�^-��>�Q���#�k+�Ma!J�麹T�F;����_=HMz�F]<0p��747V�&�dю;��vUi�ᑨ��9I���ö�i����up
���E�5�u�W�A�/znHnm�KkHÑ�S��:��Ѿ��f��S��h�mՉy�Ns��R;���V��K��]��^��N�U9�����*�}31��\C{0�z���vh��e��/y�8�F�a�\��6U�X�mT>R��=�(�1�R{��_3��c7`o�/�Z.���CU�QrcuWu�L��([z�r!�˘��'w"���U�[�Ƿ�:�m���F����ow�6��2.���3A�'2	���Ul��}V�;��$Cy�(�v,N�=�LVX|��F��_k�j�sgY.�MTnR*"�K8n�����0L�Np�eEt&
9M�O�
������徹ri�M��bf�5�vB�/�х�bu�}�ή��̭�ݴ��װӾ5�JG�u���g�v��r�a�K�.�Sכ�Gw����t:Z=\����v|3+��x�9�wG"�;���=Z{���m&�7��z�rػ��.��59�6$��r�F��.o��@[��3�5_t�ք����W���λ:ش*���g:3�:�E�qƸq��n<%!{��F�e,C����=��(^ʮn��n�	�Y����y����y�ҝ�"��}��������.�]�!��1�(���1�m1�P���w��}�	Č�E��7y38�P��+sc�+4���4�EU���.T�k9�M��WQG-P�P���=:u�[,@`L���iv���z͝} ˷�p�eۘ�=C4+3+7����y��|��6g��gq�W4�_�R8S�k*G��R��*W^TCw��%��,k=�oWM��l�5�ʡ{d;����bZ28���#�&a乓�b�D�&ٳ'v�����

���ANL�t��M�ɋZY�yMm�������+�Ӹ(΄���mU���j�3"�ċାnI6>({��v�T���z�����2�r�[�LUg��h�"L��Ӝ����\�r�KHov^ܷR�u*�Y�[�&�떺���o��̫�+��5K8kehŹ��7jS��YC(u�V�}���"�4�t;
�&�1{����6��h�����{�.��^Ep��x���T���ĭ���'&dn�1zhY�,η�c����Yng.D�{\8CI�H�+zV��QW�W)�f��U�@������k�F�ȣM˫���`aeDe�Aa�oo$h��d�gM3T��F;��wVF,�vevj��;IY$�)�tu���+e.iU�H$tK�5p{����d�j�6]/&��v���@�nkUitQq�X�*a�������}��tE��K��i�^��H���}UVֲ(N��;+P�a�P�����{ywVhZ�\�kn'�d�6vv0������zfU[�N�����I��w�d_g�M�cBT0���wcb{{a��}Z�b��m���]�ZGh"��2�:ڔ�7�����l�(s��mk{�]ַ��:j̤��79�A����w^�w��GGqVҮ�#U7�"�]ҭv7b(Sl1�F�r�Պ�V�mBa����ZZJ�)���(��V
��vY��F69�&�#!u�O�CN4��:*Т�t5�zK �T��.�`�1s�6�� +��b�6�w+o��Ӗ'��i} �w��hܵ�^��Q��_t'�õ���k�̿q���k�͔�R�:p�L���vw�e6��v�2&�-s�d%�d3������7��0�n��wJ�:�i�zZ�!�3)!��c�:���&�ѥ�l}{o�e�eV؁�U���5�tj�5ē���/��<�nTvGV�b�O8Ɏ��;��\ ǌmd��9�6+��T:(UU��$M���=U��ƅ*�]���<j����ypr��Mm�+l�=ɕ��Qy��f�Զ�!Y�1��"]Ǎc���X�C0��ђG�v:6��WUetCp8����J��{�ڭp�ʷ��벛Xi7��R_�X���t�џn]f!�\ܱ��K��v�[ܶ�k�\�I=pF�f�֮�&��&Q��i���+��p�g9�F��t��,巘��^��XW���2�}f=���e��R�ܶNu�1�W4��LUkD'�IC�]*��P�T��vC-�C����=�Vb]\!�݀��	d<T`��n�5��e�Z�+�[i�c9����w�[��D�[�T.�92��CI�'&m"ej����qe�<�Sn��{�(�5��-ڮ�o�7=+E�Ř�f�[���eL���74S���(rk껼�v�n�peZҮI/7q�:x�P2�<��2��J{/P��31��:�U�"d��c���-���{e�.��Y�����m��n�������u\�H:q�:Ӂ�\vu���=9n<�{T��v�!ݦ�f�G/a� �*�
���Df�N�gM�G�����L�j�F�n���'��w��p�2��r7:��J��Έ,�͔�Taqm�7�z��i�oR�f�A��)�ψ;��%��Ms�kc.�|�ne�1H^:�y֒�2NL�O	]d�/r�@��o2*�Hʪa�~N��y �9SV=�Od�������Q��9�����l��:�ʴ�h2�*��Y�����l�'�RQ���'7��{�.�[�:���$ϲ�+�������l�W�}�l*�Ն�P��Y���vc9�ʒ[0]��wڲuQ�栊�t�^��W]"���D�	jpۋE��.�[�LD*�''8`��ܪcE�lp̮���#�r�tҒ�ܜ�%�fu�)JpN������n�&v�P��y�ͅ�G(f��u5���ӛ��<�[�t��&[sM�e��V�j�ju[ƈK�,	�nWceR���m��Xg���U���q�J�`�UՎ��E�K��:�ɒ�s�N�zhV�:��j�U���HWZid�\/2Ge��^iIJ`"���y$D�ʒ4-Wq!Up�S�Z�Y"��^OZ��<*����jK�Vul��ma����Hx����$����th���J�@�u���[��7�y�-Ԉ���{����+��Gu��k��؋�_I����!�ƫ��Xx*�i�l�ʷ��.靉N�J����3�s)�!wmŮ��*(w���ޮolM��gq����'i���u�]��!��M��Y�uE�-n� ;��*�_��ܥN�ʧQ���nΒ�ˍ<B�8��˷F��ċ�E�����/O
��2\�FmN9�n���N`�ojmi�.!}�����̩�m�����:$�YB���u
x��,<�p�噻v���Q���\Յ�!��lm7N�rs�K��q�E�˚��xv8�W4�޽o�Ima�0��ñ�܁wx	YK��j{�[2Јѽd���.�Y�১��[bM�\qs��y���.�P�/;n<���rJ�<�&<�W��8�&γ���
�1�K�6��;�k�[^F����2�ҥ7�:�@켺����{Tol)s;
`��|�5 ��U
�.WyU��-��3T�{\fs�mg^�3j�$꫺-��;��u,��Ɍl��kZ�6Ҋ�\�O����v�o۾���v��4��Ap9qw�۾ᬆ�J��\�n
��o7��C�ZrB�m-�K3�\��S��#�C���	�kC��q�Ƴ,Ԕn\���z�L�Dr�>� g��6��u�U�*����/[<#k.�����q��������v6s��-WB��-��9Q���4�5�Wk��4��뛙���;9���*--`o��7��L<Uՠ�Ga�1-k���.�RZ���3{2��7��=~��+�5Y��*��+u^{�՝�5͗��e��a�<�Z���27��;'Ljzj�T��c��\FEI��n�>��)=��Ɉ��2lbS���fٰ?����cݶ6m�3�f���:fa�+�¨w�_����A$m��fgy� ���@g>�Nn�﹙������ޒIA1��$�F�0`��A�!���w���8u�I$�_{{m�I,�m��'���WW�Y$�KԒ�$�I%���/Cfuՙ��� �� �Ԓ���q[��E��S&�TU�T
B�nlLoL�j�y9�(#�*�!T.�]s�⤝���z�f��`�&1d�[W�vUTk��`���?X��Mwɚ��%�/z�s~�Z�]j����Q;x�;e�uomfd{W�vN��-�X/R�8�t��"���G�v�elm�b!�Y���}/d�����Cx���ڻ��{��9�c�-�n������\���¬��Na���7�n��S�m�N�B\u/�|��LN'pmL�}i�w[Fؑ fH�Ҝtΰ�����n��b�R���MLm��ݐ�pSԮM�R]�p�yj�w�zq�Z��*��a�B��6�D�����U|f���2�E�[�g5]�q<T�n��e��SJ��|�D��X�I.��N�@��3w�v�ǽj��Mu���T\������3/��^S���{��?nwJ[+���/m�تt�ܛ{�*;��i��q�4칡r�eꥎ,����եؙ�P}�D�������H�uKg9��vj�m
`�,aeK�X�x�;�Kߣ9�7����7mH�[����	s�f�/R�%z�7/3n�b��N��꼌�!�*�{Qa�u�Ug���	:l�&n*�Ji�E��(#țGX���M�Gn��$2t�Qδ4;�\��<rN���{{F�Tm�����ۄv8�	81�����//cq�U�v]��*��z�/u���J� �Q��*�NM��i�tW��RNě��^�^v�JɌ�&5Cl%�*r�ۦ%3a�q��KЂݙY)�5��V$ղ�1Zg��FA� �������]P����Kcg=�6�^�)l�r󖥁ۇD�8��u	�Lh6QUL� Q�G�u0��b�T~�x�B�-�nh�E��u�w� �e��0��A�(�N��Gq����� I�Т��&�[�v7.�je�WIu+�d��&Jy�۬�c�T(��)5B��V����m�I���
�}x��%ܣ6@4�����1(Z ��D�!y�X���YC�H!�H���q�E;�V���1�]�f�:	�Jc(��a[��q���t�˛-6��+t�N��Tl�D5-�;5��k�v��X�0Җir�
x2j�|;k�[��H�	�N�( [c���%T�y�q�Z�k�4!c����M�ݺ��Fzj��mKW�����`���R�X�7��<�-���`TO
/,w=Gp庎�����͜�}nZ���S�����[�ݞ�rW�tBa����o��/��D�@���o����ƍ���*��$�B����j��� =�9�{}�x��,E��B ��S�h��H"&�$q�L�iBMi�q��ktV���We߳0�q}$8��&S��(.J���O���s����e����)8�(D��f��!�X�|Y�j.ӕ_H��sE'� ���K�zhC�!�CAUF���j���&��}��w}���BMfI�ǐ�"IO�|_�����xI�0p�I5�A�
����z��̼�m}�����Ӯ�0:�]�� �!���6@)����~��/W���q�j��| � a��1x�n��=V�1a"�2v�U�۾F��R1��T��8X�I擮tۼ�D�n�WTi�O�y�x Q��@g�Gf��NW�uc�q�۸��ՙ׮n���W|=�J��s�o.�u�a�4@��PBEB��
B4b����[�=MUK��$U �L�9�h�+u��8��c���Q�Ŵ� v��{@ٯ}0�9��P!@����` ���!����%\��a��B��
�G�I =vA)��,¦���*���3JB#$B ��i��Ǉ@6����yS4S7� �(I���� ��0�}����|Ŋ(p"�k�@�x0,[�A�$�{�Y�a�,�)8�P���OQ����ǙH��P��X��A��C����(ot'�4���O���Ȋ��@�>�6��ڇ٬���t��?�}�7���*R��z�b4�����4��iC�Q$�9Ekn���wR�8Cv(��<�mR�d�w��]K�����q��q�5�ȳ3��t�*�[�I�7�'��g�������VuW�r��RG�$=��(���鶩�UU^aI��!�ď|��(�F�_�Ufo��������I2xq�=dI#���sF��e�k{/�s���0b���,44 с?[���![�I��&q2,�>iE�^�K�˸"
A���rC@�A�!��]{�Ͼ�K�� ��-���� ��Ax��b�+O:�{*~ DP��l�G���NWƐk5�eV)$ʚ���v��$pܲ%��<7|<8��ﴴ��X#cP�2���"5�	��~����4�(*�A!����@C�����9�҇'|��:�1{�>�����"���1��=^
�KZ$;^���s@KY���g��_	ޠꆩ��kl0ŎAy4X��$���S���m��y3��!�oKm��O#�BC�%V,�o1h��R�c�;]ٔ�|��Rt5&�N�@����T��� ,H2�"�@J�!G�E��nH��G��(.JA=G�!�S��W��\��cB$P�� ~`���q�x?�.�ə#M�  �!��p�NJa<zM��RX��58��S���
>/~u���v�&��`��]�$�����R����c�䤇$E�TǬPl���pB�����C$ar� �"��&E�}F�Y����ة�-��b���C�|�g���xm��84X1���o1xP���!��eu���r.XLYR!%r�9Z|Al�-R˟i�+x�{�l�i =+'W�����J@�n���?��b�ńV5��z�]�W�%�MjD�{��e���c��P�����̊\��ͶT��|.��Fj�:��o4�f��ڙ���1j��y�ܝʮQ�K3*�7�zF�-L��m�1��i�"���0��X| ���rޜ��,�[xrχ�� �g��X��C�{%o��s3)�B��S�c�!�L�hAX=�,n����{mf|·B�!�9B#����c�,�ɗ{c�N�ia�(Aa�Y����	�����G���0h��c�!$����1����|��w��d>����I'�
�rS���X�F����D�=c }BF����G(P�|xb�+�N]D� m�8��H�a��xI`��]�'�}��^��`-EC|PA�X����!c���;_}�R��U�ai��&	@��BHt��j��n��;J��~�C>���ܘ���H�����2>>|{d�1�}n�R�%f����қa�(8p�ƍ6��������oz�-�����:9��B�VD�V6������k�dj�T&�M�&��B�,e/I����ꀋ ��<�V����H&ߚe��6��F$|=��G�{ �D��@����4�f��V��o�]����oIy����@��>���Hʩ��EX�d�9T��4��!�<k_�2��t ���	vq�2KB#dB ���n=�$�����9V9BD͆�'��-k�������&�����w<A~�r""<�����{+>��]��� �6�,�fAIxE�bo��&/��M��v����B����FJ^�� �/�8P���GǏIb�H�h\��·�"k�᪇(P�i�xq�'�T��b�A��8��2t�Ͼ����-���a�'�k����Ц^�Tz�b�Ծ�ԟF�(�1IL�W=��T5S;!�=W�{b�[���Yr]]�Tk�'8�l��w�r�eͨv%oj����+�%�)� M_;q�5�P�9%�ӌ�0Z�� ��m4x:��������)`��QZW�����}�}�l, �4D����D��1�$��&>ɲ��~q@D�@�c��BH��5�j��r*T�#�!�D0��Jh�M����_�9a��>6�'*JD"�@�����Xo|�3ٱ��suY%96��ψ-�B�sǨ�ш4�_�/j�`�F;8���X��!e�)�{�id˿���7�f�fI����s��x�fϾ�m��h���H�D�v�
���}�rIfݝː�Aǆ�"p�
Hs�(D��Y1Z��E�\^?Ė|<�PN�#�p�Gݜn��	�߰�[��U���]��*�ә��H`�c�|��Ǆ0`}�m[�c-u���ܧZ�j�roh���1���8�(�]�����rAoanj�X�E��$�6k'Ŋi1"�.T����D��������BIQI����*e
t�y$:�)A#2� �%"좨�d��  ��i<9��Y_i��z���JsҌ��3��Y�}��4{��O�̀��P?1�1A�*�I#��N�\"F�Y�9�	 �� #�Q��@1�A�6���%!��|}B$z�I��P��d���o�^m��C8L��$,2!��.t����D�L��h��4���|A'����*��{�zӗ%�B La�!%�)��I�q�>�T�4`���E}&��%��o��}�����F�D"P�2���4C;�|Tf����{'�{!dm|�����v�X�1�A#�~(��>j��!�&̬�!�7�èֽS�::uUС��[��W2Ajs�4e��:�6m(��}��X��UK2I	Y�X&ƌ�-���8��h��eA�v8��<PH"		�H�h.�,�G��("E��o��@��ް����2L���� ��(F�F���uo���"b-)�ϊ��A��i%�Y���Ϣ.~(�^���E�1�E�}F��Va�d�������H���O�
��x���z`��^L".M��� �����ݏ�@{���h"������m(0ŉ��������+Ќ��䈑�*a���d���܇���Ti8"���"I0�DP�$Y��*[Y�[{�}y�4J�2H9 ����"Dy�،2�c�EEL� �O�i(@�g�>��^'=�,�3Ǿ��/�e�ȏ_�^'RЛ)D�"O�Tw�ZDV/3��!��I����a�M��1��WV�����1o�0��J�}o)gu�2�U;�X�v��᫄�ㅇ��1��Y(��H�TX�tB�N��ShĈ'D%R�a��"���%�(���10b,������J1ʤ�<Az��x��*z�G��UX�����h:W�~��x�2�=��;L�&�>�#X�~˄D}UL��4zcS9(G�>���8�`��b��&7<"��N�YArP�>>�K!W�~]���9��X�"c B,�|��挽��ɽ�uTjƋ�<�|e	L#�Ǥ�3��Q.�l��! �ECN�P ����s~�r6n��L�b�|�I��`�����>ݿdEM椇<"Db(���A�X��cG BG�J�_��6��3)�7S(q&��'`�a����occo���ԛ���7lej#i�<G�"W�(�����>'�$�a���ec�#���:
����\/L=S7�o��U[,�[���v����I2�$��{+~������w]�N�G1��na��ҽy���bBHi	~~���������@M��I�e��v�M�N+Ƿ�,����A��;����W�M3��7<�����"�*S���me�#=t۾���{�]K���t^��=PZ�8���,i�r!2���pW��uę���]{�7���e�M�м7�H˴)�ke[�Z�w��J{�SN��j*bͦ
h�xC�_�q+21����2{g��uJV�x��.�����u*�*M�F�n_NVnUq}��n�_j֏��Ur>�oU;��Ry�T�#����V/�^���|�ZX�DN#ywm�)�uOU���5�x����=��.�w�;�=���5ⷪ���}��!��3��Y�j[�wa���4��X"m��b!Γ��I]�2d��\k.����\�Qe,t�!2�YW�V��h���/F��{734��BY�٫kF����Ӕf78ʝ�Ah�CǇAA}ݦ�H�C��n���@��9���"I$�nI�ݒw-6	3�ř��������I$�K�-��$�[m��$��n�ܻ��yy$�K�$�]tI$�If��-��x�m��.���I$�˫m�I$�[m��$�I$�����:�b
A � ��ْ̝H��mUt��m��o(_UTT$ ��Ez�������\���N�LUڒ��+�s#G6f��i���O��u�0J�n�Į�X�51�&K�W�f�DT7.v[����k���ƒgk:q91���҅�l@�t5�O]HM�Z�J�x���{Y�Os��Y��M�R�v��y��Ӹ����;dO�{'H9Ӓ7F!�K�f���G<wZ��ٲ�Je��pr�|��֍Ӛ�rƍ�;����:� ���ӓ��ûDU�)����Fi��V����c+3�rΔ��D�`�A�N��8�ju'[AI;_\̎]��(W%��I�5���f�*�2������To�Յ*�n�.j�f��)vs�����:侗l���e�g4ݷ�5-��77�G�Y�M����YP�W����۝��d��*Y���Ow�mrs�>��-���,��[�Hr��wz�S��yCc�S�d��A�S׹/�q��HδB�ݢ�>��pt�p�-E�{���$;�M�3R{�.���J�Uh�>X��[v��Os��l�We	�y��ٛ�+HA�ʢ"�HT��⪱Y|��Ղq�gHɧ	"R0�	�ځz��h �H�%`7:�"U1�*O5PR]�]⍹�c���ue���#���e	^��]@�Zf�8;z+E��Iф�~�eI~��J]T�W��+#j,��73^���]��&���"���L:�p�U�T2�C�v��dV1F$:�|�n��B�e��c��C]ЌPjWb���*�D�gt�Q&���/�e����5�ô� ק��*�ݍ7��9��Pe�2��O<`ķ� �D���e�p>��4���b�J=u�I��e!bZ��6���A=6�x`�W�,�yUKJ��P��f]���OS��Ҙ�b�R�2�Xw[�Dw�S׻b��<�㐼���On��r=lm1-�PA�";l�����4&K��Z�F>|����`P�V�\4�����0�6�LFX�msA�ˋEQ=�Vv�h:<tZ�[	�_V_M�yU35a��;�/y���x! �@ �AZ.ΫH�%j�� �*�vt���Ƭ����k�j���g.����T\JοZ��J7�H��DP6F&."�/���a���vtM<2i^�|�33F��-8�>}���=���ql�3��:p�{M�='��f��?[{�Dfu<'�������@�	=�8�[;L�è����8�ۂ�8�l@8�$wL�Y�o��n�~|�������t�r}sř&t�S|v��?-����ˍЙ��٭�8H��C�	}�ϴ�wu뾟X���2���^���~OI���[o<��#x���]�bd!����k�
�虙�l&�2�<p�Y��Ǥ�3|���Km�뙳�,�f?Q�z[{[l�,@ ���x���%�ٓ ��m��t�ݞ�gH��^�!�G�>��#KoKc�2Bd&4Cz�4A�3Ĕ}���TND@��d �09���!�$p�c�:X�f�ù�ӎ�8t��g1�0�f����H���n�~����I�zY�C�2Ghv��߾9�����ϟ؁3In�: s���υ�}*l��5�[qś��e�����&��sǎa��,����Hz�<!���I��j3w>��3��LQ��̖��{���9�ǋn�$ǟ�3����-�}G���!���L̆c=����E�-/<3����L;H��V����9"�Q�1}��Fc�P���[W{ ��q;PPAC� ���+�J5^e��1�+���X�W�{�y&�˖\���`)ENr�å�vٶK����t�KɜI
l����@�D����"b��^������<A�8��n[���-��9�����{p�d��G�fqm�[�xLxD�n>�'�TS���c�3�3��&���,�1b��8΁�&	��N^}�\��^_�8fq|��4�!����z[=�8�Kc������g�:������'���>�yk�!�o�d���Ä�p��1�m��Z]8�g�߉�l��&PÈdc��"�q��nfs���;믯y�����M����~��!�n�ߖ�Yۜ�i�������5	����K>>�{{��6��&􄟫zv��vn�����&��<��s�t�Lv�虹������j���5�L���|8�&ryzO7��<�&��|[�䍸�,7�m����n�}�C�2�����Ϳ��O\�u�Kt�g���#��q<[m�[v�}9���v��C:#F�_{�j者�}�p�0�>8�gK	�[m&Z~	�z�
��F&fs�0��=������v}��!��Y#�L`��h�A��Ә�ӎ�zGi�X�
��C#D�&�W������S�֣n� χ�!���h/=�y�+E���N��5������4/����]�c�'��XuK���8XG��)�t1av��\m�kfm�}Û����H鬕�I>m�(��m�\��J_U��|/5t��2�U�͑�a#D��Ui�I��X����t�|�������y=���i�o~8�{qݳ��>8:Go8D8xMb�� 8��ߥBS��M�?|p�8�����,{�-���t��x�V���z��왙m�q�����-�9�D9�nV�4�y�q�[z�Ӌ�~^���ť�[uӇ�{H棙��ś���v�cy�B�3i�Jڳ����8��-�C��d`��Y�uBË����陙p"�j�y4�69ɰL�#�:��ӏźOHqfqx�ٍc'�>���QU�V�ȱB%<�&���z[n,v�W�zq��&�g�n'��mY�����-��9����3>�}�g�i3�2P9#�=��9�{M���6�w����H�g�C.���AP4���o������oI����Yۜ��>'�yzq�x��ig�9zz��6�xB�n$~��Ɇ���I�x��\]�kM<q�d�fd��hvC��P���ww핯|�+�� @W�� @�#徻q�K^&n-�X���~	��f��u_���5/}�ft��K}��g�|~�^��ex|a7�"8�D��3�ч�~�;"�>��X�)-���0�0��aa�Ul�&�q�U�,�r�M�����7��k�6��`��k�U!y|�Ǣ��_cT��#{G,zK�#��Mڳ�ؚ0!��ڷw`4	�O842 A�G�����6n-�O��Ëqۏ��33@��Jf���� �7������̑�a��"��~��6|N��=�q��3�q39��O����v+��g������:Xqf}�}9����n#�m��m��z��Zǵ��������$��sެ���<̇���%��	�q}�����#D��*8�7�I��>NQ�|St��U�0�ԬD�
I�M)�qÀ[�z}Z��f>8����q�S�B"q�$�8��s����ק?�WV�Ft	#t��P�d@�I�}=bc���" �(��jIS9�:",wM2��#���r{.$�(��I�<�(�7�X�z�3i�V;�řd�Q(Z���I��9c���k#��+��LL�&q�
O�C1ْF8�D1C�O��	H��ѤI\�a��˾V'��͋��I�,Ě���m�Og��PX~~��hD�՚��(��:����Q?G���)@����%����uѝI˳G�+�c��|�#;uη�6���vά.��>�GUq���d}~��C���b4�)����#6)]�{o�V��� Pax}�˷9��=/�Ǟ�m�Xu0H L0��I�,��W��q�%�`a*��/`���$gkbD4&p����>�)���F�Wo����3"�}�X!0�|Y>� {a�@��v�bY36`�B���	Fy�ޒ��8�����2�fq��lC@�eT�
L�W�pC%�vK�Ǔ̼�Q�Θ���tC7p����q�>'���
�0�7�{�]�E��cxbcɂ��g_&gUI�:Y��Ǉ��,�M�nfv�a����W�VՇx��`u�;c�����u�{\^!�=-��B6G`a��RX����Q�2��>3�֜�y31�R$`)X���+��w��877�{��p4u���=U�}�;�q�f⎩�M�M�cS��3�?]��ű}�,�fiBC�Y<�}�����~Ww7�ca�3��b>�d��X�}v&�iDM'g�������F�D�G�!� ^-)���i*-#�wP�eQY���I>��}�-T�U�T7�o��a�> �A: �ܙ�gM3F��"�kr���y�n*iN����*I�n!w�UV���5o�1<0�+M�'.�ᲝfdO2P�IH��#�~��4E�vu��Jz<<�z�:�?��N)���a,�Dh�=,����X�@�B�N�g_�c����Rh5K��9�h�jv ��%"t�F��g���0��?��#nD�k3�����Q��$k�I�L��헪V|�!s1E�ƺ�|
���2H�c��#��6����,���D���>G
ɉa�c��C,#�:�Y3}��
�v��OT���g�mn�|���2���g�>� uT��+�\T'G3��{�O�bOq�X�Ic�R8�ڱ�L�i�!�&s�W��t�TC3�L�|� G���s)�wR9';{u���������z�c��K�'��"!�=VS�f(�f���<���xD}�مTUy��qz����/|t�#����d+���uI��rڤ";Ԧ�[����O��)m��4�K�n9��J�	�<�F�^�Ll�^�u��vBXjV�!��;A��uUL��7�vFS�;A3
%�ޫ2�ž�2G�������:O�{Y.:}4��v�)/;��p��H�A?R��b㈪� ��)8��c�uݰy�>��z���8��`�֙��}�ļH͒���=�BV\QTa2"OT`�C�&�d�Q뿦=2�fd,דҕ��9c��:4�:��q.�Y���껿01k,�h��8���<G��r�u��;�Y�=w��V�3+���<w��N��4	x��rV|�Yh�%ہ"��ǘ���t���d`�C��U�l=ڈ,���!=�qԳ�[꩟31�X�F��Y/aS����8=�:$��{ߥv�_^fS�!*F�FW�B��p�>��[3?0��RW\��Ḁ�p�?�Q�ߒ&�?mr�g�VUS��œ����P��9��*���@�T����hѣF�W3AS�9��Z�y-��}q;7��9c�͂�Q7��[�r�I��Ȫ�'���M@�ue�wkKd�hR
n��	+��X�1�L��B���zc�K����8���r}B%�r�����Ì&]�=i�>����t�D�V��
JH��4}�e�j��3��w�D#O���1D��"���3=�4ۻ�ɴ31�w�:	�4��ݬp���d'i�e ������٢j�a��d�5����q �f,�a�R�ٙ���@a��`���
3i9uCu�38��4;3J Cq�=8(X'A2����s�CB�3}�vOn����8TD6�ď'�!�	�|m�9Q&!|�~�u�۴�uU��V���N�0��΀M�<i�+qْF;�A<�Ii����@���h�1�r�a�;��!|qt�9����U����]��0hD�~��m��s�ubȌE�
���ҝ��i:��X9e)p����/8�	���5F�ׯ��#�{�@ߗ�zO��n�ͪ܅Qd#�89D����M�5cb�W(��Q��� n�]9�����IvP*'"�S]ktÆ�g#�[u��7,UE��;x]�6C�����4�a
��ց'&8&n�"%�}������f�1��L�P���4�}��:��튼EDAU`�C�N����}o������{��>/^d�
�t㎣G�K�{p�U���2������q�'���y�.K�'�z�i���}~���Z�����G$����/��RDi.P��i9�����1"��!]Yy��
����%�w�gDq��]n���0,N	����s�M�-�$C@a;_��������4���28��lE�	0�\x���~f���C�1c��� �������e&��X��
������9 ��C�����B�`Ѭ�1u�EJ�<K�(� 3�׈Y?8��]i�;���`�"�~ޛ�v��^���9��H��bv-��7���a�3A/ ��1;��J
;b�T�ۘ�U���w�]��۵�r�CL�:���kə��W<jdE ^�D5�1fMA hS�A�S:��s�q�?�
���!C�$�*�(r	�v\��^z>r*T����-�(O��;?�.�VC�pqY��_�q�`i�׎�Y�"��L�c���Є}\	�f�G{j��i:��Af')d:���'l���I��{�˨����>� �Ǫ�{!�'�B'�J+Y�|aǉ�t
�������>�]����'��"8��w؋��́o��"\�(On�J'��*lwሿv���w{�9,a�qW��%��JH�%����2�|�L�L��C�(�J��*j�y��q/bn`��}�Ѣڬ�65�pC��e;$�h'k��_��������ըg�#�~i�:��gFrT*��\��m3J��9���B���ӥ��x�:��;}�i�vW��>J|��r�Iĝm贳c��Ӽ��+Y�ܻN^�o#��%�^�i�]V��ml��;m��v��8[��W����x��r���T����l���7X"s+��u�
K5�=-	YW��gm���c*�ӣ�nφ����Q�-��=�^�/f�n�u'��w���y�yr�C{���]���=�����ƛ������V�
/���B��t��k��>Վ�y�[Ձ�߾1Я�A����:.�r6Ѹ�[�y��c߽S���E�:נں>�q$l���[���NX�o:����J_0�A�Y����Re���i�2��v/i_��2΋�e�f��,�E�ϼ�u�Ӈ��_!Q���|0���eV}h/`uiG���je�11e6y8cmj�]۳+��ӝgMw�Mŧ;�ԙ�%�b^:���O��뵑_r�Z=~�]p�y��ǗV	}�K�C1��t����
pe����=J�i�ĶYG�U<Uh�u�6�����U.k�=Wm_ʲ�r:���#�W��wK+
n�]A��2)�v~�W�pv�L��;�TEs��Dת�5xۻ�?�I �	0p9����<����}��l�{���I$��&ۉ$��ERK��wݗk��o���e�Y$�wu���}��=���d�I%�~��m�Ie�m�I/����]]�d�I/RK$�I$���[l�u#y�������I�ղJm����.�u�(�.Z;���iĩ��Zfw:Xr�n��k�s�,U8Ru٠�IΔ]x;�#Z9^���CZd��Fq75v!z��{,miJ������ZgQ8���L�ar���FU�:4o���V��6pcm����V��M�m����r�u.��tt�u�#�k�*G�.جj镼�fGl��er�"ts�qR�� ��2Q�W2�w2�%�=$xv"�4�S_j�z�g8�l��ٔ%�0ڳt�=��+���jL���r�<�#w�3s3u�ƶi�X�z�J̡l'FVzH���7F���J�sz��.Kf�Z����qs�n�]'p�I���%jԕi n3���f��sZlE-)�7��bD�����p�V���Ī!��W�c�Ƶ��k"��m-��EL��jF�5� �Ǆ��F�mu�䄚����d�0X��-��l7�������0�ƅH,���sS��ٮ��\kV��;{��j�[��bH�Ÿ�s���M��Tj�e2w���w��*���Y���f��Z�x
��鑾">N�9o �|R�b��q����c�[�4��E$U�~~�=C�fދ�:%�����WU���fY�ê�t�ۮ�{�r ��
�<9�s��$��3��]e	-Z�.[���ku�aɞR�ޢe<j�)4��|��������}�w��6�H,�%Fn�q�1�Bt�j�E�Z�I�'�!&�S���o��JM˫́%P�ќ\��ɳ%��ݮM�C�j��4/�ѽ[����8��%���v�,���z��U��U�5E�v��T"�hT��8'ղگ�o7T��;0%�E��ԯ�f�2V�Ͳ�[qc�[���a��I\�B[׌N�FhL�2�Ao�m�*b �.�0jJyT��U7M1x��Sm{:R��Jq�+cmۢЏ;pۭt���BFD�]�Q������oS�r�s��bO)�A�P)V�)��UC�	/΃�$�3(&�jA�P�y�Sq7 �Wan�3(P�O3TB��P�9;��7��~#��
�iV�AEq��tׁ�]A
�:SE���qU�/��P<�HZ�ȭR��y&`��<ޫ�R-�)��v�NC�4�ne�ٵ�|h� �l�m��R�P���%��CZ}�۹7���c�_b=�lE�	0��u�K�`����>�D�8��!�w�I�Ĺ��
ˊ*�&I6����n}�35�{GrO��d?������,Oc�}Eu�����}w�3x;��r�F)�J1:��	>���~���"G ��0'�y��8�D��@a�}f�3g�E�H/������lA��a@�� ��)�}�>�mi��>��4|�J0�z��C�g���г��r ᣶Ϸ���xM��.��\.�� ����	Y���asͿ_�<F,Ac�X��/�	��8�U��>��siQ���;{_�!�*��	��ʖ�!���I~ä5T_�,���~��WXW[.�x�H����yCD3�,�^q M@�%	��e������.�-�~���xhѣGx0���Cq'P�XV�Z޻]s(��������8Ry٧jU��1���̌�D�VU��D[N��h�&ܩb����ZܱY�`b	�\�����+J
-�PH��0mh�� �E��n������CX�ch�C��&,Mdd?0nM��O��8�❒D4���츉uO��g�_�gE�����=��؅Sc�M<N��7���^��}��X�?%��	��U?T���W��'M��~OVC��R�㉂��;��|8�e���<�Ew}���Q�#�懡��x��Z5"
�x}�h��ߧ���̱ˤv�(�t��&��I�������၍���k�D~h�U��=ژ,�I�಻�<}���4Rk�g≻)�{��r �8>1��� �C����P�K�� 9�3d����ʝg����y]ڔ8�hU��l���ɟ��xҊh �����72��-ٔ]��u�{;&:�LwMO_o_I�,���R[��f��Ʒ��cYskXV]m��X��Dn$���A�A$��!�@�#B*�l�+��ۙ�wp�?QF!L�tFa��<L0�w�<w��DG��=�]&\�L�9������_hB&	c���r�Dv/[��	��*lw�ܓ㉲��ѣ
��e����:�>P�	�wF�<mY션������rM��A!��ğpj���G`��Ƣ ����p��J&!��s��#��r�츉uO��}`���}��r:n��,� ��B���D�'k|瀄ǽ��G���"������}c²⊣I�Ob�U��!������	ZcA{P_����b{�@>=ge���"�����ςЃ)x����"
Ġ���w���9;���Wt儠4B��w^��Z�@Y�<���U ����f���,P�זU��A����p�pB�
v��_P�n�T.�O*9{r��inF�[ɺ;%�!d�$���8^��@�eZ!h�@��ZjD�8X@�@�B7hU�.�5���Nv�oh�G���������VZ&	v�}�ϴ�&*lj=���B6������g����8�B��"&P��YK����(��8�Nd:$�]^��{2e��!㰇ER�¼K��wA��خ�����>Ͽ:s~�h�V�����W%��ˁ~�6t���u�2����Iǉ��/󼔑�}��o_J�*�#��>�ԇ�U��Y� ���Mk1Fn��wq�|�}��X��y�,��5�������Ք�a���(������I��g��%�aK����8�չ�e�ع���X_9B0��u`kR�!���ο���/布�>�A<|=G�Ć~@����S�df��
4V. QDZA�+�|˳���_m6�-���]�!xh�#��R�[iXu���]�4�c-��X�ɻ-JI����Ć�nP���:��_j]�1��@�e��O"J1z�� �g�yt���q����vT���+1γ��Gx!?1�|3v�!����V��x�7�˛E�A�K�'��4᧬�I�$}�xh8�|蘉�2��8�B%�뼎�ǉ�u���0�����&n��5NY�+<�*�D�.�<�����oݛUJ����� �B/ʨ�0h�2�V/����>·f`�`�T�D=�?@�3S_{�o�ns.�-�BC�J�]�C��G��l�L��>/=�oi�Io�B���*�E�X@��*PI�i����=Q1A��w4��vx"��W�|"
�<:�_��p_#�VMp��A%a�
�{H|�F8Y�ۛv~o������/"*�Ə��+)�Pؐ?$"�6�����݋��XA|bCC&��U�%����­����F1e��2J�:B�F]B��Nʬ�ɹZ%[�%ۭZX�mAC��#Ȃy��%l��%�}�x�S��1���1W+��n�W�%#V+G����u����.�#Z	��b}�f�|t]��齧��]��9���Sc�v�$O+Da���X�����"c²�5�+�3��I�S]�[ٲI1��#����E=Y��R��%��=����g�/����;��}0�ˤ�i�G��'i�pQ>7�"��g�G!�	��Gm#㉲l�H��=z	��s�Oa앞Qe�`�kHtx}���4�n�ms�yu�+��La�r��C�o��\�,~`D�{��;��eDLP�C����!�T���pWx����¡��c�Yt�c�28��oh�}1�ڒl�±ɼ:O�Y�"����������9kޛ��i��)q�.ל��F�8��cۗ�,f��kz��$���%���9�ѯ��l�:�D�%����"E����.��P})1���E I��/���H�q��7St+`�E%�HD<S��y+HČ�]^wam�st�*���XC�R60@�2(w��.�=��{//qD�¼%�w��#Ir��;�G�i��D�31���,�B�QQǇ*i�y!��^���-߽>�Z����:��LP���O�a��Ȯ�������u�D�x!�OX��"�� ��k|i�$N��7��%!>z"�&l[t)p�A1�ĜN��OU-�w>,�OVC�x�)�����G������U0�:K=��H��#���vR;Ƒ���O5��5$y�뼎�Gd��@a��p����,]j��"`�kHtp�����;꾉կ����<*�g(�`��Is�����������p�Y�o���Ƽ�_;����*Q7/���$�i��E��2�,]���ۻX���K(彥**��6�d��dy�C���Q��n�*��^�Z�	ε=����^�8�A��Ia2Z�gв�#� J#'̂C'�A��q��efl�
e��7
�0h�:�V/����v:*G"a���ߣ�������=���Ơ���tU(�4^%�p
�<�ĵ�vth�q�]&Z�L�9�=VC����]�u�}��S��=�<%T��
��b�x�<q<7�n�r�_dMXag|K뼔�K�'��Ha4m�1^�X?"K��[c��JVM���k#!��:���������9�8;:G4��3�q괈%�=����o
��O�gx�L�V>�Q0A����?a���Woe�.���\��E<x�I��}f�����bϛ�;S֐��EO�r��;��ц����~d���ƾЎF �|>�G�|N��H�Uy����L���+�V���8��N��̂}S�
��R<.�/O6�(lݮ$ף�D�JǷ����_Q�٦��r��Grw��O��8� 	�C����U��*�<|�g"����>$��m���Y��d��_V]��0�59X�')�H�A��	�l&����HۅQ-dvy(�l�!�hO�VN�?��ƺK15x�D�c���P�L��J`������a��Ui�
�A�Ĺ�<X�E$A������q�,����s�c|�J*LĻ*�p��`��O2���I�]�X�L�9�>�!�w�!PL��D�3U�,焧�	'��	��w0�����/�ݹ;�a�ٟ}�Zca)��BzЭ�<Mv[7c������:��4h��T�x��&�2JgsM&y���m/;���	�"�I��g��%�|D�}��.����	�;�eJ�H�~�K������о�!���A����?a?���]���lg��a�Y���)躭e�W�.8HV*��>u*�:��n��a���g+E��M�q�N�q�M5�����Yɳ��	f˔* ��(`��(
2B!�K�#)30`}�[�����@�p!&*]$,P�J��y�0z}<}����^$.S<��xV\E�L��#��M����X��d�� ��A���)XH���8�.��'U�ξ����׏��N��'��$E��yh�~����ř_�n,�4O�4M�0-jP�L��g�y1}5P�@h�C�at!4>�R�>(��E=��K:����5���0�/G��EIA�3C��4�zS�a����7wX��E#k�]��4�.��⌿f�Au#�c`A
j�V��#>L��hÌ&]�֜��8�f�x�>8�4�
�RH�1���-�2;ru���/����1]v"ׯ:��лV��_��}]����z��3��*/�R�{���xN��^�#�bw[gՖ�v,h�fft�����^_(�?/�A�����@�.��ϏhU+"���>�hesI�r����w�N�B��`5�c"(����Ajw��n}�7�}��ʥ~y����i�6|���m��H�{uOm-ow��=�鲦$+I�)�7�mWR�V�����ٱ�=�:�����Xឹ] 5;�3�ŻX�����TZ�����}��m�ٓ��/�*+뼴_j[��Ȟ?z���Vpf��k#�h�o}d�w3�/F�S�j������E��w����{�����̤������1?Z���ޏ��޳�����l�����ߥf�_�}�RZ����k+Β��-�g&{���g��D�mз��eVw9�b_3�|�	|���>�d��)��fͷ��֯1�%����7}��6*����6d�����Ô�M�8+���_:�,e�E.z���9�θ�w����.��*+dרnl^Zިdzg�_�����7��s����|y�5}n��F�����}�/��`v�u��/��!���EP�*�Q�73� �-���s�O�׾�i�]m"A a� �/����H���3��@C�#�������>���8�fn�8e�����ww�����$�I%˖�l�Km��d�K��������I$�~~r��,�I$����-��y��m�Y�ݖY$�Kn[m�I$��m��$�I%�����.�%����$���RNH$�*JNqR�9fUk���`~�����/�����N�<gd������z3����;�H�˕���4��\�gtL��~}�m�}[Ns�WwV��ewd#�����ZIBFv#w���Zv+���Ȫ�K2vM�[e�;//!��1`�H�5�om��$���	J\��v��ݛ���E+��}�Κ"����=����Gl������yN���V����2Y,T@�Uyz�θ̴"�}.���9��s:�f�ڌn:��'��!(��s]ʓU9|4�PmŮ���kƮ��]�8�5�=D`O��ι;j�w�i�ļuW����*� qSn���M�
��g6��<��j�P�K9"7��8�FRQyyA�褲U��ǆ9��s�j�7ޭ\�IN/t8�5�U7O�v������5����}��uIƲv�;�k�.L��Μ���s��Mw>��wY�[k�AТ�/^��˗���-�͢-�3M��Q[�kv�'R[Fgd�ig9g8_E�M�n����R���Q�2�/��n��5H��nīy1
�֞�'0h��3���d/NGr��3�۬9�����U�s2���8\.�&���v�7Z��<6Q�1ܩ
�R�7�m{�Y�~Ҋ�n�6p��3�Pj�5���B�e��fN���V0S��l�;�\p.w+�sVI\C���͗�ҩ�f"U)Z�[շ�U�����ƮӻmN����A	#NRu��]��P陭8�θ:��ͫ����1_nY�2�|BJ�%���(͍"T�A#��kZ40o�eQ'Is�w�Q]��!l�L����O���^�|�ݚAG��lh�שm��:�Hc�.�ĴZ
�i7�V&�R��AR0!v�	�2����Z�5Tv�K�򶕭��{AW[N�1ErJh�)t����{V��H8ro=ʣf%3ąW�w�kZEE�-��a�,�n�A��h��(P��˖E��h~g�b�\ܗ����#T���o��˫y[#��q@�
�guKǶ��/f9ms��Y풺��I��]ڎּ�+���mV�9	
1����e);-��D����J����!�$���EN�4�"D���@U2�aQhVek�וj
O#�L���U��:4u!�ї
�DGǇ*i�0f�>�m��F[�&m�<�Kؚ��u)��i1C��1U黎�z��������{."]W�+s���aFm'1�i���x{�� s����y��>%��x�>��;&�u�yy0dA�[Ga(8u�)U��/����GS�fҎ"�s�;��zˤ�iȓD9<Ay��B`;��üa�H�C�H�M�p}�gj���������	���<NQ����&�D�#�Ip_���2�k�a���ൊ��P��S�� �A-�l���q�t���(��&
�7�5�C؜��^���ɣ�NG���θ�>?���4kˌ�̳�������uTҥ}î�E��������7A���/ ��c����{��n��F�v3��j��m�۔j܏;,A*��\�����*�W�����h�p����L��TQA4�/)�"K�>,�e!"
�(��nʜ�ʪW��s�,@�E�i�l�#����V�������`$~g�r�!��|j	 �^���Q�7��_zjj(� ��χv��&�,�\�ܒ�9�Hj�i9����i�1Bq-
&�Y�Q4a�ʚ�$�4h$�Of��~��hd��D��6�d8�2��`��ěZ	�8�����a��0���rL�%ս�I���b*K�4�7���X��\I�W�a`�L��$��H���������ϳ�I1>�ha�#�B���X"�H����D�����}�}�F���h$��.�w&�>������>9*q�CP����D��9���q�l��rv���AjU&K�~8��� ��{��,3˼�
��&�I��u`��3���
k����[����ڂ]���l�)�ۼ�R];f��wT͎�.&dnQ�uurꮡpΣXEI]�vj��j��2�Y���.!	rC���I�TAed3!>��/S
��[�m:��c��$���v��p����r�CP��4sZ�`��g��w��곒IAB�+�YF*({�w��H6ǂ����߳�˨��&ȣ��D���A>��N*�h۾0��˺>BIL�Y2<;�4r�>��L�y&Y�<I�p�W�;�F�ן}�2I&$r^��QpJ�9B9��}��*���$�I�H��I8�
,F�	H�9B#G9�/��$�)E�HI��BB2�Ob��N�&9P�8�lG3|a>���mV_��B�D�>B�(����0�+��f��a����OuU�HBHH�d�h�"��x����rdvs��>�c�ȏ�2I!!΂�h����+�TWA�'s�j���2o���/�YK��?T5��������rL�K�>��F%�m���WR��/~��mk1�F�a��J���������om=����8�e3K�2����ON݉���㢸�wv���%8�B6��^�d��*���$A�,p��f}̐�!��	�x�RP�"I4�'���M�vw?���@~ֵi��������oSź��!�IB$Dxә���<虉�&I��I�Fb$�H$È,D����l��ϴE}.��L	0Z/LC�QC�">Ơs,s�y�O|h���ϟY���fd��ڎ>0y(C�Zx�����NA�f��<����kL$̐	���Ř��,r�9Tx�H��o��lؘ;X�u�X���g��P��QͥE�^�3$	0�1�l$� *�I� r�8�4�Qd�;~��Dp�&I�Ŏh�D��(r�G���G�9�uQ��d��N���(D�<A�d��68�ۼ�M�A����oȼ�� i H�g�6����Ѱ�T���U��ꩱ��dh��ذ�l���;ٖ��K�&Gk=��i.a���8�޼��*�����z'��mvq�.��׈�۶3�cfA{S	D�5�Ha�<}q2M@�P"H%PB(�O/*b�����mʅ9�#�!�4sJ�hIZ��ܪ��$��������w�}�p��,�ȡ�.�Ab6d�sǍ��prf�{�s�ˬ�3�ZO�XcX��a �BŊ"3a�+�"I��9��!Ib5I�Ğ,r�9Îf]�7�=tE�{�ϸ�sQ�$�C�%���AD��>>��LLDy�S$%��	 ��X�#6J�d�(���D�XԆo���OH��Ϛ�̱ɔ��4y8j'�����=Dxi�A���rI� �Ô#�{�������3M���zK�ʤ�Q�� Ev���ꯘkI30"+Ė#��g��(E�i0�e��	��iw�j����/���E��ʂk���/�"8�M�����#�P�Н��z�!c�Y��8 �$��ޕER��n�d�v]�T���swe�&��F^(u��9��q�o,�JT�oY2#Fd��R��%E�/gr���,��&��)~��n��>(�(C���Qb8
�v�������I��Y�E�QC�"0qHx��Rv�3�W��=0�f6�<9xD�� ���DJ��g��%�m�fH��c�L��9e�UK�I,Я������t�U�1�.>>�X�L��q�d�"9���0��wd�Es3}ɴ�L�"ʢ���&��hB�����}����`���8�N,r�9�Ǭ���^xE�T@���^�!˒�H���A�HI&�k1����os�~��������H,D���d�VA��)A㆗����*#�R#D�sP9�92���㇒�fR�n��Z)?���fO�(5���~#�@}�z|�Sy�Yd#�/�]O��G���]m�~��g{:h�8J��A�[��N�Hmet����x����_H�>�
Y�ٗ)�����Ҽ]<)���*f�.�6�s#���XDq��6E�C��99�j�Fz?;ʸ(�b�pWIG����Ϝ�i� ��"osa�]�Җ�fOQ$��Rr��Đ"�;`�m�p�$i�������s��P�i0���U��$E��+�� r�8�<Q�#�i3���Ҭ�����F)�YAT��O�D�^�;wK�|ʣIQX� �D�i��(s���g�Q1Uɬ �;��-ʪX"HdGxѺ�#~�.������2C9㏤�"!&�d1<}�{ޅ��fe�o�a{J ��l4�SIB1�{��������8��X� C�i�$�X�$�fa׵=B&��W�w{0N��>�xQ丁��D�iVF���X�|����7��*U|ԯ��Pϕ7�nX��A@��|��Ĥ�n��s�i7˰+&�mZOj�&ߧ�=g:��b�&��F�e��q��MH݋�Vsx�����3J�N�Qy��0
�bb�u"#w_�PD|Y���	$��� �
#�����|����(L�eYdDIHr�rDs1��پ�Lʙ�<c`9�92����%q �f���LY���5�&���(D����>�����'��Z��}�r���HEv�ώ6�,Fp6����ٙ�t}��zLB#搃(��T�Q����_�|�&k��6�Q�ȂR<A��]z�e@�9�ÊÌ���;a4xC�B F�Q㏳{��������\�$��5(qϏQC�������0�wZx���|"HE9ÏX�,F^�/�ll��3�zPǯ�(y�|؟+1�$��۵
M}��>��W�u���3��$񤄴@A�*en�ƈ5R�թ5s	ֳ&�A�#k\�{�e��3�U��7��K�}5�9;`�T�ng^	�l�-��$��D�^�6�
%�$'U%���$�����A`� �A����es���פҩ���� �D	��M%�I'x�y���{���|��N F�sL>��E��M��B8k(��Sa��@���	$sJ>8��H�z{>�jYuw;��q�R�����si۾�֝�]M���v��<<�8��m�Y�Q&��uN��2`� �&ÚCd��*������ �3A�"�;"�0�(�$�8�'0A���v+������|�UT�	0��#����ެ���y��8��|�%#H=C�"��_EߐC៻"O/f6����D�����rӥ�<�c�|~R�u�g�"�Eez����:_5����n�A,A��(tP��$�ro=4w��ʵ �*�i�U��v�뵈�'U8���_v>�.eZ�����(�$��V��0;�i"j�	��YT�X$C���N��:w**�N���``�?�;i%�P�iع�n���_.|Ͼ�����DrsK ��cI�9\d�l��Շd]Mz�xD�� rg�X�,FL��i��x�I-��,q�����)U'� �F ��αT�R4�bo�1���NI�(�,G��>>'��D�2	�,�R,M`�=%���p>�kߐ�
M�hI#�Q�Ė"D�Xi�6�a���($�Q�C�]H�Gj2�5��]��3G����2�6�<`�8���� ��j ә�6k�~�&��X��P��C�.�*�C��#]7��Ҵ�G�WX�S �����/�Ћ�\oL^�t��R�<*�
;3�b�F�,�v7{��y�J�P�Hk�j}_vw՛T~�3^_Gm�j��ݙ��Gj�sC��Y��E�y��G��e��������l��|}%�J���%�G���ɜ�1@[�8�߽'v�<��^��<.6/�mwg0u��zn��;�ʃ��Ej�ؾ'��s�B��_^�Բ�Kk~c�s��u��g�����s�p�����,g�8\�	pfC7��ɥL��Y�]�[�<���T_
:��e�ɰ$f�A]�'־�D��CM�%Ѫ��m�*�Ч:]�+���K)���mڶ�g��_,��zSײS�=�9��Թ@�)v�n�`�[x�N�Ov8��P};
d]
�����_l\�ڱ���⤾;��.�}x�2�隺/���wZ(��5���K�M�(n�I������8���M�w%~�c�UX�|Oo����[֤�[��1Mٙ�X�4|�<��>�\��Q������f%�o2���xU��*��X��ʯ�U��I��WQ�8!�ܪAw)y)Kp9p8{�9B�^��2Gbۻg��*[��U��&���=|��ٟ
t��D�k��RLƩ�����\�kJ�r�3t�V�s-^3=߮���s,�$�����3 �^���u�wtn�����}��s��~]^^I$��3:���-��e�Ye�I$���譧;;�� �&0`A�ö�$�^��l�[ן��{��r�$�Ԓ�$�I%�� �J�đ!�kvKa�A$IAw=y+��b�R���F��t.���B.[O'.���tP�jEˣm+|0M�g��ⱼ�wE��ʌ�#���7�*�7�Xk��'y��$��L�+����!BBW:�{�w�����q-��*��n5�ĩc˼wy�ܺu���nm�`�U�۽�Ec����f�n�<������]�A=�wVRҦ�u��n�9��X#mt�\���Y.���_<e�x�H�9	��MM'�
�{^��{�#83`̝Fw0�>.�V΢�cs��f�Z����&b�Z�a�ٝ�:�͢�"`�z�h	t���!2�mlT����S�N�q��ȟu�Nn�r�o��k}Ɍ� ��Q7s��}��c�fx�V]Y�#�q���v���M��)�q�g���#Q��w�ڹj�����,e������]r��tx���s��1�gLb��Ʋ����[��q�7����S������:�5c���y�w<@���}ڙ�e���w�Fz�NPm�Y�
��|kXYJ�c.��l}{�&�^�4/p���{MN�a[ٸ�"����K"�n���-l��TYѝݓL]��ש,�V̺��/n�ۼX�n	�6�Du���ʺNd�/i�nĞ�6��(�.u���P���Diă��U��˪�p��]*��dyB��yJ&V�&T�a����\U*��P��s�d����B"]T�U8��v̽V�3(�W{�����P�B�.>v�(��[�2�%cJ�&i涅������hr�OKH���N��:�r�f�y�]*�ŗhCx)�i<��V�#�A�<s-9�̣����F��o���������݅^m"��F�Y��fd�^qK��(�h/��<�v�u����Ej,�a�O������32ߵ,I&{���Ε�/u��Υ�cqӔ;]�)�a9f�MU�����j��2��T=�3����(Cڦ��T�{�e*y�nI�^A/"�j�Q����'�^��2疍����ka�MCb��`"`*�	X
h�"����#T��ML7ء8���GC��<�*��1,�
T��n�9*�����+A1u�;]ϧ:괂�tXc�7��i��!�9���_�K��,����4[�J�&�F��E���<�3tt��4�U催N-��D�������h��>���2��N{�?��2�,F�0�9�P���V���U�f[�����
�PI�ÐP�a�fÈ'�lr�_\M[Z\|#Q�Y���)+U4��>&]ݙ���k,�%����Y#�":����뻿3�x�0��s9����U�UR�G3_�rs��*��|�a���ȑ�1���lI�i��g��z���8�Ǝx���)U� r�A�Q_rrb>`��9��ߓ��qG�<�$!��G�=�qG�~9/���5A�"D�%�s$�"0�M�I��o��HۅQ 6�9Q�"D�^4�e�b>�Ό�j@F�~u��٫�k��!����K�+�Hz����a4�O�����U��[;R��{I�P!R^��<4h�ѣ�EC-�nZ��dr���Nb��Ƈ[js���K�i�6��ь^��C^q�[�r	��˨&OE��>��HZ��Q�T�`���l�I��OC�gΥ��&��9�`䈋����N�(���ֲ�ݪ6.��^8���,��&��P�f��;��㊻��`>9���=%��Rr��Đ���}X+�S̼c��N�K�L3�|zJB#�B��r�N���`��	�(�P�aǊ䨱�+}s��]ٟ}�Z�0�� ��c�C�j�QBm9��w��ׅ�e�������b�DJ��nm2��xF&�rN��r�r���$�Q���ݮ�_:�횎Øcq�Ȓ�i�H�p�=?�������f�$�~�
E�EaD9B M�㚚G��$}Խ�E��=���߶j��ϔ��X�u�_>"Ћ��Ԡ�i��<�9U䫏�GT�E��ee!�>m�8X�(!�%���T��|�7wt��]��ˢs�vN����AwvΑ�kS�[:����b�C���e��!���R+tY�Hi�)���ب!�`��+��$2G��	4���1"HC�����G;~���l�ް�o��d�"DG��
�,��OkE���V����?���D"d+>>��Y"$�9���m_�:��LA�0rځͱɔ��GB�`�o_���\� a���	� �\�i� �r�H�M8����g{f�F�8��NUi$"�;`�ƛd��ė^��Au,�>E�;�Q��"�G�!Q���8�e��֞ϋ8C�!��|qZ�#�i]��oƋ����x���!�Q(�6|"�ѯ��{��qw��<q��br�r%sI4��/I9ⶹ��.�TF�'���������/Y���f/O���g�+��H]Uv��&CD0�cE�a���9c�i�7�\���@����G�V�G����5��o.�餥V=f\��;� +��}I�QE�M�v�O�v}8���?Z�U�_�\�)���}�4TaʱʪZ"HE9�N���ȅ麰>��֜��⏎��G s>��s7�q�d�n������qd|f�A�"�><��V'�:��ҥ;΁�Qg�$!�񧬢�bh�D9��9Zy��Bf��8��0�Se�I�|q��]�]ϛ��y󍆜&B��A��A�D�� �H�1u�|O��虉��F�l3Ó)��<�8���l���qՉ!$�� �nI4�p��7�4��}c����ﲼ�v]���!�����!�Üx�$��`�ߌ7y��D�Np��$$�C��'�P�Ɛ�(�
�ZIF���5w��s6�CC�_;�s4�-�?w�W;�<|��l��@҈ǵ�K���Nov�,˞��8/����[��*A%�ET��`��*�+K����f��;La�V,���H��y��Z�}�H�w��W^�X{�'y$���7�a�$�� f��]U&P�R4�H9F�9M�ME@��$\���%�(�d�ٮ8��I'ğ�}c����,GȂR<A��$���^[Ѿd�	;i PQFQ(�6xE�B F��AǏ�]n�T��	 I�(�Oi�L�|I�"��a�s�y��f�����!�ʣ`�r8s��/�s6�}f�%�Y$� �!��N2����z�-V���~���,�����? j7Đ@��&���M&X�$�Q��c3�V�n���� ��!<�}e�D�s�P�f��ώDʜ`���6�!$�Qǈ,D���p����d�Ǵà�4�ȉ)A�(����j8�g��w�b��;YFB�Xi��,~VM#�S�|O�U?:�>�b7���F ä|}�,(���il�ԑh�"��w�k��%x^{Yv�!��0�6hʰ���ٻ���	���%����N�-�㌛���E�ۻ[u)�&��
���h�]R]��z��
D�A�%.r�U�/ڇ����$D
����>������~�]Q�!Ӂ��]=��P؃pB�M����X�Rr������U>�q��X�D��9���c#���؍����N F�HAT\�+(�C�#��}�g��\\3Y��N/EE��A)A��F�p͕��f��4�~%&�NrP�8�K���}�Ѣڪ�a�H�s�0��@��s��9\�������]�T{�Z"HE9����H���w���E0�w�I���Ah���(�4bN3���1�UW�1�	��榓�8I'x�ȱ��gg�ݟfUd3�G��E��M礡"<i���'�m^w���m��%�}*L�鸄�P�s��|p�Ou�{��������Å��(P�7��ǮU�x������Э/��t�.��]���uՕ���{�+w]-���ɪ��Zm��K�4��оD�%�m!HF`����yv!J�X$B�R�h/#T.[��B-�����UV^�Yj���	i�iv���f&A�MVpI&�Q��X�!a�`�9�����>��Ƙ���9���|�e�k1��t�Ƌ�>��ق>Z�q����� ����NA���Fo�ੋ�a�,G��SHd�c�R�,��G|����c��s�:�,GȒ]�8��"�k�������ͻ��2@�L���A(����r�8�4�mCa�e�?G�s�̡T�jD�߿\~'��R<A%�B �(0��s�GU:��ҥjT�*�"��IUi$�i*�����;MƖ#$�"8�����M���}��]��|"V�)��Z�i�֊KV��,��$���"��x�M�ʱʪZ"H9����\��g�o��#�	'�� �� �kQ-�T�T�շ�N:�����/S�#��(�+�w�N;���}�v�m�#퀤ЭJ>ע�ûΤs�}�Ѕ���6� ���m���w�w��+�{��M���b��B�!���$��F
ڱt�i����L�oKs������L�w#ƅ_KV��y����H��SA,-�^�UR%PN͚��[Mӥ@�[	��/�R�������$������[ZCıh.ĒV1j�5m�����>�IUQd�U�n>;����xAh���(�(D���]'L�X�	L�r�o�M��I>(�"�Iq��v<����}����30�8�H�$�C�%���M�I�7y>��Ǧ&�ĎA�x��H�6��1�Gn:� ��C��99�P9�92��qf�Nb��<|}�OQ��H��*��9$ӐA���͕�^���]�wH�<����QXY�Ev�f�������Kɤ�#Ǥ�!��r�>'���C�GX3i~1W�`�(C���ƖQb9�	�v������>H�	)�a��}0P�L��ⳍ^��'�^���v.��֫@ɧlg��Z]��L�����ԑ�)����>��lrX��g9�17tUÔ�{.	�_U�u�Ujg8�[M`�^��kKQ'�����7y��n96D�ug6���o�vW�@�n[�"D0|�@�L��.�*�k� Z%�O[�Qj�CRH3p]�� �u�����a)&/S�	dQ�DK�2a��`�q�"0�,r�92�9�G�9���*S�M�̈́��qir]�]�UR�B(���8���Nt��\��؇D6_��#��Q�h,D����$��wd�EX��㈿�5U&�A�7���sb���D�N��g���>(�X�!���F�y���S$OX�y���B$D|a��$$��4ϖ��{�{���ك�qb$L����Z��R���b�\��s����Y�����re;i�g
B�`+O�D��37�³�'��Ϝ�* �
"os|���O�+���dX��G���+<P���M6�=����}�!K�+�������`Ջ����L��"5a��ۊρ�>����|�	9ۻ�,!\,0�.1��e��:��8�� ke4zeʪ���;GGK5������ˠ���#E�rȆb!WK-��6I*��KA�q�O�(����|	�!�a�,�lC^tǧS��>֎�Q"�]�
Ộ��m��ϸqh�(@�y2�A(�>2�~�"$Vq�ABMgYE�p�R8���ͼ��U�U�P��C��|AG�
|I�&�e���J�w7�ŜP��,���re9�$����|}D�TH�c@⣤������!@�#�s��ܓ.�������r$vs�z��IXA�j����Ͻ�B��32��G�� �&�O54�c�3{��������i�qh�C�>z�-&�4C���o�;�B2� T�d��9�G$Ѩ�����1�&l(��VQp}e�y%!�>E9��v�_�}�\�v�ͧ��n�Ls׫�ԝs�Mf��ĥ�-L�fu�B���yR���>�����*Sԏ;<�t�ֲ�3G_111���r�.*�����9^`�����3�����z���\�!��d��XD�i�N���wI�.�fa>d�jz���w���}%�ke���:)	��ʡr���K�)O�f�}�~����1��Jg7�^�ѿ5�XK{H����j��_f��Y���q"ܿ<���{;:*.��+�304�Ǧ��qH2�֋��Ү���:��D��\�]PU�UZҹz9�ezn��|}~^�ʐK�	,�x>EK�zB��#�]Rw�[���U�C֟K3��z�`�ss������I���"y_w!8���ޗ����2'����\x�������i��u1&tw�v	�{�w6��i��j�2�yޔ�ԿF}n�#���_����iHz^�������XU]2�W�q�(.2��>���8��Ո}9���q!.��%�>�ϯ}]��(wu�T��U�S^�g�#S7�l�wWׯT��Н��uҶJ��³x��$�2R%��u�<5Z6�D�_e\�΄X����ͥ��U*�yPn�&K��l1���� � Ø��o�y�}�� @t�7wd�D��{���Ic���wbѡ��w���ﷶ�_I$�I.\��d�[m��$�_m՜��3��˩$�K��������$�\��9r�m���m�Is���,�I%���m�I$��m��$�I.ffs�\uyygwwrI-�g�����~����f�۳��v���I�dOWW]^W#۪�eԳb�Ht��S)Ӗ�̑�B�$��Χ<0;�:ol�V��:(�ʻB�xQ��K)��Io����P�(m�u�4�i^���/%.�
J��t+�v+���gP�Ud�������
)fF;QuԈ�ݸ���\�coS�I�v�q�pS�W7>�+"�*^ԧY$n�tyݥF�p�
ܤ�?�Ϊ���8�Hlh^�{ z/ql��U��{f��[l&%�W<]|^�wNwS��HU)�uh��l���;#�$��걁nۚ�ɽ+c�ysJZ��Wz��;�@��iF���&5WW����|H��a�*q�9Vl���O0+d㓯�U}����J�稣Xu]�iW^ȕ�8�,��=���=Ɔ�@ڙLp�T��n� ܮ���D��r���J&����0��DS��bJ,.�Ds��Q~T)�NnS}}D��#5�Ua�D���Ѝ��T��l���.�Sy��a�4r6R�N^&�aV�����.lV��<|p�����Ţ�uUSϏLuX�2�$L�UdW��5s60欠�age,
Y�b�������Z�E���-�d�|�z�Fm�3���s(���J�]�[��i�[m%Y���X�se+Tlu�����ޚ�qH8ͨ�ՠ��E�6CrFU^��UK+׆W��Z�\(u�i�-���C��p\�4�̶�ʎ���]WH*�La����՚���6�/���E�K)�w���׊�dv�4h�V����b��ﱋ�t1o�x^���!|���VЪ�n�h���Ӽ��	���WWG��\G:A�B��&Q"c����()��2S����9�]79ͤŞ��B��U�<�"�M�ܸЭ�GJ�ݷ�6��Ut���.��6C/����ESQ+RK]b|�����U��ڏ��I���~��oՔ1n�:���'�s6�r�f��3��B�$B>qCk:r4��`�n�Yz�� a�\ס����}��T�+����B�d����叐"&*�D;���Y��f.2
�CF�Â�,Xm6nV=�[�	��;���[�X��6��s�m��"��ޭ���{e��,�Q桯*Ůt��P뱄3�8��1�a&�N���1z�Tj��'F����!��|O��'����*�fϙ5a�k�竲�Hd~�a���re;a���8����������x��\�* ���H���A�5�xZ��>�]�S��B!D �di���E����a�y��{�ffe�!Q��>g �>�QE9�#��w��eO�D�x�&��H��RJG�(����oҶ^���OC�@����(M��rP���8�7�z�������,s�NL�|Q�"�8��8���a�T��9�R�D��ak �Np�u��ff\��g8���B�}^PZ,�f������iEu��fA��5�>ji2��qF�o�>��y�N��Dc��a�֐�1h~E9����!:�IoȌ?#�W�x�3�XѕA�f��A�hAC�����t�&֣��,�ޮڕw9�m���Y7��QQT
����r���y%S���Er�Q��H؀Q����/!B�P'ʱ��|�Ȁn���F��'�Q@���^%��!.}lsm���D����Qh�4I��(Ge�~�*cC�I�
�쐒M ���,D	���^�Ͻ�]]�$�Ì��8�ȉ)A�(����������mi}Ou<O�A�j,���A�d#�(�Ov��|�=�$r�(D�;a����J(��q=��]Ua�� q�b�s�:�,F&�P�$�4�,�����7wW�& G�c9Q�J(� ����|a7��N[�y�Hq5�Q�/��HI)AG��F�A�U��$���c�O#�o��7xE�B Dq�X�3F�ޟu���Ͼ_l�Ib�9sJ,��@���0�3]��R���ѐ�>���C�/��P�#����9��E� �>Y���u�~�{�
��t]屌�]�"�,`|-.��M�l�v'}������\���V�wٙ
Kd���i��=Sr%��r��Hx��Chz�]	�cM Ϭ�f��H���)Q	�gJi��1$l���2����E�8�Į��87n<C����$Xs*W�I�E�|kY�r$vsN[��X��S&L��>��B]r��eQ^(�5�/|�OU|��&Ba&mbo�1���"E�(�,G3Y>3��{��TL�	$̐$08�q��Qh�4I���"DF�A�x���~C�|�2HL��HI%qg�"�Xi�+W3��j�gC0�$3%b9�P��$r<9�s,�5��U��3G����I���6�x�HP�O�>��X�����9��f��k.��B�&d�HBHa�P��4Iv9(�����n�[O2��ꢴ���TU}No�߯vIz��%���(G���.ǩ]���I$�I!	�&,�g �2	E�cP�E�?!n�����x��L���f�;Rfi�%1�8��*Z���'��5'�}��e�[LS���]�s��o� �0�0��X��eĤ��Fl������:,�Owmr�BIao3}�W�>p\�|�P�{��,eJ'6�aI"Ty� �н��]�)�e��XG��Ɖ�U��$�C!�#4�[U�d�4pI��ݴ��z&I&Ig�ڨ$�� �ܡG� | �x'�Y2��42@�I�)Yg�(D�� �c���jCD����K�w~o&B&M�C�ad"�8����˱ʪZ"H���N{ݥW�ϙ|0��2G�x� ��/S�#��Q��sz�z�,��d�$��Q�^ ���ʢ�QP�hQE}�Ɉ��Ĝ��f�"�y"HC���Oo�~9*˻Z�2%r9ȑ4Ib�(D��4�Se�s�o��J��*u�M�AEAb L��OAZ����Q:yԻ��HrE�8�a4�e����g
N ����ףb��á$�&�G� ���M�x��o=�2� ��F��r�s}W~��LJ���E8y4���>��*^x�#�B l�ƂTuA0*{��s��|HI�r���:��G^�3���P��bw�j�zwOd�Wf=���gU���֩Ok(������S=D���Er�4�Pp�WL��wT�m�q�k�z4M�R�5�-�-e�n���m�ᢼ�����rQEag�!ۙ��~�<���8�v^'bIB>(��8qA�m<��15��+9�"�����q6x���N�mj��b��3�W0騄�x�(Dd>�Q�	�ዱz������u��ň�,D�> ��/�(C�Q��O�/>�`Ħdxv��'I�9v9UK�B(G����ݮ�_����&c���n �ND��x�M��B8bȧ��~/��I@�@��4P�}d�*� r�@���54���G�D��5 Ha! �>�aĖc�"C��u�f��\��n��5	0�}gs$�">> T�d���c=g�3Δ��������`����!��J��W������>#nC��#M�͟S�q%�7��$�A�G���;`�	=���6�+V���M�5q�v2����5�	ϗ�N۽�ņ�c���
�q䴫 �k���Q4�m�&Џ*�����E������s��x	`��&B��l�EM �}���&n�Βd�KJr0��G6�"Go�,�(��o_���\�6�L/�M��ښ	��G�Ӂ�	�z�ث��Ԑ��&	��EŚP��9��'&o�3�{��O�BBB��g�E}AB �� |�d�S�{�0�w��&BB��8C�igH��7�5��G��i�wk�$Np�#�?�]ABl$�Eɣ5�{�v����1�h��� ��/S�(C�Q�5�w�$L<���qi2_�.�*�p�!"�p}ſ��1k�9�'"Gg8��
�!a޲	�>����7�`6�=s>n=�k�;�D3��}(y�C���xǡc9$b�o����l��g�:P����ѰҧQ'�Wt7v���Bsd���ɷ6�g:؁}G��s��;��N�Pǌ�һ²A	���ـ�0$�*]݉�7���%'3��D�����HC�O�,P@��x�SI�8s7�u}�Jw����$���BQ�-&�Z!͓��N3R��G�{ T�d��H>,�f>��������>��G	���p}e�y4��9"8������3�Q� �H�xr$v��g
B�Xi��2,N�S#��MiD�;|kA��X�0}�^�+Ηeݿ��96i�Ev��6�/��Wa��t��ʞHB4���0r�6JE�h�f�徿D���	#�5�Y�+/�!$�x��9�si�-�����Di �肌�(M��rP���c�� ��C)| w[r,��}�}�D �����X���+b��]�|A�P���)3�'�~aۋG�عc�� ���UO��Awz�1��agwFy���Ҫ܋k��g�3U�V�RJ��\�%��u"i�Q\�W[��)OI�R�Ig�c�sn4/r�e6�����.�?��8!�'&P�>(���qa�p|Vi���لǏ�s�ʥb$�P�#�>9���9��F�����;9e��� �E��w�~�~��/�{���1'� �?�6>ji2��i��w�=�n��ffv}:�<By,��-&�_s�P���>9*m�FŒ)�$�H�qg�,D	�����/<W�ɿ!a�m� �T�"�rD9A�#��o��=���wUY�	ee��ag�!C�,4��dc�q���*S����<@H�/I��R(�9��>(�UQ�	�#�p�!�k�� ��(~�A:���gXn��#-L�/���DC�Z����3j����w��&|��WK���A�#�!B���:܍^')<�3�vh�ڝ�X��;�8]MR�w��bY]���f�169k�8;-��H��y\�BWs�hEeF��ygfY���GΰU�ɣI)�23�9��F��)�ŒBC��tr�.JE�|!��<���U^���A�m(��Z^�	%#H(�"�8_<�0��	0��h��(M��"�"<q�9�|a>�h����jf����aD�,6OX���o����ۺ���#�J�B(D�k �ND��xә��O����8xD��]�Z,�(�rN3���1�SW�h�h>>ji>��D��Ės�#�>��3���f끼[�>�}e��iT���H�#ƒp�Տ�}�D�O����HD��YĖ"�Xx�+S�1h��wq���*���rD9x���,r>�6�.����9g|@{�0��,m���z��@|E�ڀ�Mr�!�qg*���J��#���1�H!��}%�8FI��]�Q��m1��k�wo'e[�5�������i7�����j���T�I�$L*NB&m�7�t�)	����or�4^��3�0��"i0҅!C�/}� ���9�J&6�3}�L]hň<8��+�,r�Eag:9��������F2,����;J�������>���F�ŕC�<ْR(�0�� �&Í6N��4߹�1���Ґ�R> ��P�!�, ����s�GU3�q�\�9|AŎ^'8m���m�J����� Ӊ
 v����6�.�*�h�#�YFo��Ｓ���}��d#QQ���^�"Gg<x�h9�g<���럈Mb0�+ ��E����AB M�3e}�uU�"�o�M��D��Ėy�8��ǘCߣ��fYN&���?M�^ɽjো�BI��D�[F�p��]	YȪ������T�b?���X�����Ѣ���geJ��F�pV�\�@����Fm7�e�Ձ2��~��+���:k班��2N�ܵcF۪/��.��םwge7U'q���]z`�թ}g���y��ub�sc��o���Ƿ�6����k��oW^�M�[�-��My�sF���G짖h��{��K�oe:9^x��oL�G�<wژ�u�7�bZ.�Q8K��/���]V�j?vO����{�^��e5"oa륏����|iU���o��~������)�o̪�,�"M��j��ݐ1Ԛ[��Z��+��ݷ�{F���5��_5��k�B�A��b�����7�ͣ|�ym`�ٲ�PY���H��.��O�n>G>)���,��U�<�Sb�V�{wa��O��Y�+=un�����~ܶ��{�o�<�qS���C;r�K�Wf���Խ��\^S׳�#Y�}b��}X|�i�RH�T��J�^R�:�(Iw<yk!TU8��w7��/�mn��N]�UksU�QY��+�O�P�5f�t���٭ؼ))�Cyx�nӤq��neũV�bz�����6ܳ2�H��n�9�^y烳�"{�fc�{��w~׾��s� n���������I$�w3:���� ���Ax$�bnwww^�m�ܲ�,�K�=��[$�/om�I?w�����,�I$�����I$�K���m����<Ί�Mn�ѣC �$�T
Cp$��PG� ��r��F��U�
�cΛQ�kS��")���Lw����ձ�E�kB{AT���p�3r���T�[�ܕM�7ԅ��:�[z�W;��~J��\�k@ƺG���C}�[9���1�)��Fd��l����{�v��\�a>^?q���0�2[����b)2��ڧ�)�޺���[��i���J��s�[����Ƥiʿ�(�yCԾ��Wی�6�P.���Lj��y���wj�{{�i'[M�(���=���ų.}�9
/�Z�Yx���y���yl��8z�ΰi��Txh�+4U�g{^\��˥���e�2�բ]�1ctb'Ke=��f�ACۏ��ޕu<�)u�Z�l0�vqvr�bS�^j�:��ȣ�.f�31r��n<I�l��T�)ڍ����u�(S�ޞ�����ٍ��YY��o�)j�wA���]*v��=��F`���Hj4�WT{2�<7�����; \�|�J����tEws�c�p]���g��T����"j�QJ��sr]���!�0��rf�p�����z��{�NҐHCs�8��{B���X]U��	z�pw�8I@=U�'����Yg\Y�N�#�����n�M���Nv�}U�v�.��4݌rvPx|�vNaJ�J���	>UL�*��ɧ�+�}�5t�1�����x)�,���ޡ���HbN�ڭ�4�Ɔ#k�Kq�Ü�- ӸVb��Pz�բ#��v�|����f�t)���w��b�$�������w,�{�H�[]��͕���A4Lyq!�a1�d�Ƕ��୬'_�[n�`i��c[7fN]J�e���Vʘ�㒫+�Y�Ң��	��tvh��i6D�&jJ*�RX)��(r�TC�-y.��>�R�a�o�l򇞕�u��p�[���kc8���q,%�j�:���
��*���d0�0e�BR{eR�.��!��g'���h���X���#!��iv�DW�n�!Z[�����x�S�"�$AceJ�Ŀ/P���I:���`�s���6�o����㖷��yX��ǥ��Pqa��,6���q��bGB�B�p<[f4�Q�[*L��*Rh�b�*����U��A����c�|�y`��t�I+���/��\�k�^
S�U�i:�^enXA]�{K2��$�����D��*�"�!���"��O���x���y��0B$w �X�!a��Z��NWgn:��z�_�$C���A�9;x����Q=������#܊$qqDvAg���9�{����˺��d`���
��QXY�EvG3G���t<D�q?}�ؒP��:��A9��^�)ES��Ls�9�F��8�l���'3~�ۉw�}��bEQ�(D�/Q�ABm9�����v��b<<��9q9x��C�|x�N#��D�����ۇ�%����U.$"�{;��/<��f��5c�^�� �-W�E����d��X��J���;9*9{���܁B��c=��������1��4n��8��[��[�#Jʧ�:6��9S�s��e��2���=�_SB��hqv����ڳ��N-�;�n!&i-t��3e��͛!����15��}�&¡�h�Aa�x)��śAb �s7�a�8��d�Ewh��E��Z��3�<kD�1�/>[L��>�|?Ig9b �8�x�*-מ}޵2D�����ȹ(D�r>0�NY$"G��,�o{��=�3��D@�L6X��r��m�s5M�_�q�~0EDH�������!G0V�'>�����gga�9SA�Q#��4��k0�����K���LtC�c��+<P��9��d�3I�ok�ۿ�	���G���G� |��R4��:d�<a�9BMg"��HI)AI�՛|Bt~��V.���#���S�"����4oɅ��7u�����q6�ğD�-�Pf�YjΥ �`dh�P�Xa ie��z�#Ϊ���PVG1nk&�WsǊ>���Ue�e<+w ��9U�m�\��[����K/�E�B���#�(�6��j�J�"
D#d�A�T����>�XK[���pX�� ��	���.C���>߻t�Ws{d�L�AŎ_��(C�x��f^�|eUQ�c�*:N�˱ʪ_�B � ��3*��~�.���S���H��,������f��c�n����˾,� �P�(D	��O4I�9�����~wt��q�O��B|<W*(�cJ���8	 �~u*:p�!̢���D?�Y��;O����1�&o�MBdYE���_��4�����پ��Q8A��ͱɑ�,�(qņ�o0lߺ y���,�=49�D�qq��O�r�����P��(��ڏ�ă�:|�CJ:���>��
�-2 	���X���5�i֒ȁ��c[�[������/`�Ã1�K�Yܘj�n���/[lݔ���r��\�m���Eݭ�,r���WZn`���Ga�^�a���� R#��
ā����\v�OɌ`VǸ��x�8�!D E{�d����0���v�Q�̬�>B(��
|9�IH�����ݐ����~,E��Ï�V^�	%#�
9��z��[/Zx����
2��6xE�Q���x�ﷻ�����G�9��&P�0��
v�ņ��G�7���}3G>�_�B � ��d�������͟	�(è,D����Z,� �>����f�e��q����I��I�9���K7�������223D"�C����E�x�L�Ib5�����<��Î}'K�vL>�|Y�&�2(��;x�H��+�i�;��^A\�ghL����j�a�mC�?A��=��Wا�����Y�(vI��,V��� i��_Qz���u�7��**�壻Ji�N[�9,4�Ū��q؈�oq�6��J�-�ɷ�/f��$���)D"4>D�/�I���ї�����.�	Yc��5��4 ��P�C��$Ns1���ﶶ�EM���X�FxR8��H7l��s���+��;�x>��	�È���R(��m�$���4�:,C�q�Y%�v$�#�=G'�>/����W�w�q<gÐ=Q���+(��(G0}��{�e=g�k8��_�R4��9B� �����D���ɇ�7�P��<"�(���H4��`�߽>��ϙ��?�ڊ��K8�YC��8������2{a�z��.j�3��i"��>9��NZ$Ni�ͦR_:~���b �+ ��E����Q�^����y�3V��O�Tt��<2��� g;8��?B�6�`�A� V堰�kw	��^_��B��!'��
f��U�ŷb��&�L=��.���N݇}��.���ޙX��L0��^�},��\�x�e0������^E���]4R)����u20٩��i�&����%ӄU6Ae9��5?UqBm>,Ɖ6�!?�$�\��d���]�ت&`�<�_�[��RdzK"�4�xoSo�q�'�`�=qg�&�20��:�9�9^���5X:nĜ����r<A�D�X��x�o���'�����6�x�HP�O�>��Y�T�@���~��I9w~�8���m�R(�,�C��:ly�f&��-�s2�/S�$�u�c����_�/<%fH�:d��+(�C�!��x�d��J/�lr��{��b�3T���D���x��
7��Q2�*G��Y�=!DG�x���C��^_C�Zþ�������u#J�T$w3{Uz|����"�L@�#������)1w�~��1^̑Q�G�()��
-���K�,�i�=U[tL�Uǰk���)��35������P����3��eɫK��s/�@y#������6$ġ�.jQAH$M�
�>��D"HB>���zum
7ww�Ǜ<Q�;h���W��c���i�/�99�v�__>g xG�A$�c9z��H��K6���U��YW3"�B�e�QnW�,�"�h5Wܜ��i8��$�B$~>$���	!�4�2��};��u���Ч�K�eRdd�"D9i$��g1�����R��>f�8�AEAbh#ƞ�ls1'+���P���t�H�"�8�9�92;iG
`ʻ�>���uy��a���VY�9SA�(���ώ��8�������&/I��R(�,�C�M��3͋;�$cqY&�v$�#�PP�#� |��}�r����z�ӄ�o�n�/z�`�K�LY��`�zr��ܑ)p���Մ/�|��Mw�����ҼAh��CP�C�a�%kss�������-8��#v���o9�����$�`��.4�����)����kv��dC{JՎY՝uź�vv�Õu=N�Z��w^z�=/'�^��w�z����B>�B��>��#�s�3����0MQ��&�Ǎ�Yx��1ַ��V������W:G�/Ô!ȲH(ڂ��s����WOw��"�,�ȃ��0E�%�sOA���}�{b#!�v��'IX��Y_i�z<�'>�u���To��I0���NZ$Nx�͠�B8bȧ��~/{�!I�}dc���Zd	����)9�7">�&f��>D�gY�"!$9�W+.NbkV_��ڻ����2.M"���%��&	�sNO����}����ω �ȣ��Nf$�M ��9����}T˨0�� �D������Ş��ߖk��$��yuuYpH�8���m~�>��a{k �!�R|Α�k�-�l���p����gA�5wdL#� ����ڼ2we�_Xj�X��:��y���,��h�ލM�j\��ފ���b�8ݥ���Ad �,�,��B4|!��!���D? �%!�D��	�I�|י��CЀH��@�P��B	i)d�溶��6�M���M|Q"Zi3n�핾�˻�wr�r�EYf�:(C�|i�I�q���{��Je�v(�#��((C����l���ĜY2�l=dp�(C��ÏH��RB%���y�GN�h���@�!���]ABl>(.C����}�����!7�Lq%��W��i��p��W�$�)�D�8��=��E���j�"q�0|a�[�^�� yI�M#�YgXX����� �o���U�U��k�
!����!@@�ώ<B�,rQ�����)�~<WIg9b"q�A^V\��Rdl�����JV!�?k��_o�������q�
�Wn¼��ߥⴒ�l�1��ϚU����jc��a��80�paa�ut����\�]�F���:sWY$�jH��[�n��^�<.��B���:���QT�y(L:���}�>v����b���(�� �|�xB͐) ��&߬��q{̋���p��YQ�8��9�0�]̲`����f�pI�_y_s�}��}��	��6�������$�M ��$G3]qQ��tL���� ��A�L��|Y��i���Jt�07H�r��HH�ώ_I��h����Ӈ�}wo�1Mx��B��e���b�_��o�&�/�a�t#K�AB���F�H��ҍ�-�z%L�30�#�5�a�+/�$"Y�z�4i9�����01<k� TAFT&���Q��i%i��]���fcǋ ����C�Y!C��8��8>+3λ&>`` �$�̲�4�c�����b�<�Q�"t����Oo3x�t�%�K���Ecג���͞��q[��_N��t���ݺ��Э؋�M^ݪH�����w�݊4\����v���������.���j���z���\�`�gf*�O{gn���uR~�l��r�8�w+ۏ����v���=�'{2wG�7��(��e�w�o"��֗��W���8ݯ�E��kUO\��U
�|r��:�.vBz�j�h鷇��^�H����9sv���bR�k�m����pRD6��U�r�L<pwk5=���{�&eL�;gO��~Re��^+��k>>��R���;���?v=���cZe�D���"Xb�-��z����=��u����%�f����v-s�rwwTo�vY]ŷλ��s�\-н�[��R;�jJ=�0�h%���U3��gf����NI'+���l�vn�Q�4���`�Lܭ��i�i���s�|�P��7|:����X�j�:���S��/O��f]	r�2T[l}.��t/��(k�����*��}$����[�VˌZȣDg�VVK��[����k��\=�ܿP�~�&�x����%�I�1���[�:��ǳ��6�ꔜm,���U���=䱞�o2���=z�T�`��5��)�[���ǈ�߆ƫ~��U6R�bg�	���ZV�o�dAb�o �$���~���y���{�;;��맾�����}�9�p��sd��CL˪ˊH�bAAI$�����$��m��$��]\�;λ�yy$�~I$�嘗��I$��ߵ˖�l��m��%�^^Yd�I%���m�I$�[m��$�I$�w�.����Yd��g7w�;���ů�$(�2;�x�$� �$7:���T�2�!�l �G0���;*�A1K0-����p�r�$��!t���Uڡ���P�:�lJLVD��	ُ���V�=xhܾj�ڪn�h�c�E�ݪ6ki�]"n�<���%8銎kJ�n�(8�������ZOVu�1��+��]!	%Dѵ)���d6�qwe��f趭�7�n�u�1<{�T�;��n9v3W)2�W����6�A%�C�q�t�Ku���J{��}�aь��AN�1̓��t�ƹ��	�u�R�'4���0�M������gqu��m�կ!�"&�:�⵹��2��ɑ��R�:�[��:.�;��ӭQ�ܱ1o���cv� M<����\Jy[��*˖�/sB��Ս���'c$aʎث�U�7�'sрễ�K^�9jy��mŦ��۵/��oo���fRR�q1�[��,�]mn���фPuY2�J��^����u:l�T��M��})ٶ��-�L�]��F�S����;n���֞S�w�`�ͪ=�e qo�������ʮ����\t����sX�F�̂�k�%��p�K+��l>x�Xvg�����P�I[3��Y�o� ^���a�+$!�^�T�H�ҺѸNݺ�Ѻ��׎aUD,�T<�Ζa�a�G�D�7vţ�nUB���i3�-�<Q�YW�z�Ev����]�m(�-1w�(�bN;jc�t���R[ȧW��K{�O�gtڝ���7��eyh��PMb���X��4l�m�!w�}y�V��W]�5�Z���I��$�,Rt���K������A��#f��AO	�v�ӥUw�udJ�ܐEe4T{H2)I']Z��UYzD����0�M�=j���^�B��L�1�j#2�s(�G�ֆUB
�wJ��@�e��3D*�8)n�f'[!S�K)�hమro�-��[h�δ�8�3(�rf�%e	����&rPXdp�j;�<�Ц"­���i5LS�ͨq�b�.ȹ�rv��NlvJD�p[��-���Rڡ�����\65$���n6<n�`{Yq�/�hc ���
$��wT��7�:�m[�<3��ͷ�ґ�:ռ�8{�t;9�˵�7A�m��̛r���	�MYIh,2���%�@$x�����H4����D�n�m�<�ik�}QPC�0����9�e���In���#N}�����K���}�fbO!�9g����J$}4���1��v>�3+;��fa��I�$�
�Yr�I��,F��g���m�`�GI.��0H�|qg�,Mda��?wй��{�� l1����IʚA�9"�<x�A��0��ت��`c�r�v��<)
톐n���Go�B*co&WDs&s�����)W�v�n*��� �:<!�Q��Qx��%��Q��O}��m�fW3�I�9�%"�s
>�a�W{�>���m<Q�ЯT�g4�lr�9i{�7+�"�_��]��WW�]�k�r���\e7��r5�P�<{=H��>+ٹ�W#�EP�ˮN��0A�a�Ƌ�,]��ږ�'��u�����+n�f���6ը�c�Jvmk��6*�U�k^B�3�Ʀ#��4�A�����*�a��ሶ�'�47.4-+9�LĿ�h���&�J��@��ƒh�o�3���뻿���N}��Yd�;|8��(�[����~>�nI�S��)�D|q��9i�sƜ����
y����<"!$i]�YnWYhE�k1��W}�\vUU�c�A��?�A(�����r�q	�������뙺�oZHsM���,iT���H�#ƒO1�����D�O�y�A#�q��L�<l�c���+%�}�
5ʿ �$�<I�s�P^ v�?����r~? ��v��޲1ʚӂ_l�4�>D	��Gɖ9H������7ߧ�ŵv����~�9����>�}��Z�N��&�c�Zw]���`���*�U����~����qc���(P@�сp2��T-����͡�(����l����0(tNiЛK��IUk��X�9���%U���7F� �:�~�1."R��O�,�a�
�e2(�0��clA`��k���c�T��1-�s=d��rH9���#�(�1�q��n�4��r�2JE�,�&�4�9�
(�}�#Y��A��s�X�r<A��o���:�����1&���@���xE�r�����{Jl��9'd�9��(�,�+J��?0��������|��b�dIe���妑�<Y�6l��(������	"�/���r�r�B,��7�3e}�uU��YDH����,�"!$9�s0�e_��ϝ����5��T,|U&E�b$C���Iw2�f�#�y{c癈�b#�x���&Fl�c�c�ߺ�Q[�"-}�x^�r��$ �+�Vv�@g�}
 l�0�I�"$�&x�i�hW�RhS
����h� �/��a�B�se��澩0_N�}��3uSɗ�����(D�1�fu!uK�59���I��nU�+Ķ���'���Y1���I� ��b`�U ����ºPV��%�I%"Uy @/Q�!k���� � �/G	"�0�9���if�N��<|}���:�$�B%��
� ��T�@� 8l����ͪ*���	$3�����r]�R(�,�C��;`�3�ݞw"q�'
+S��A�:KB�@��|W��U4��	2@���#J��(C����B�Pp��}~����ۻ�?��B��A�a��
>�Rƚw�.���v��b<�
C\�D�,�Kz��d9���9�#��D�30�d3�iRQnYnWi�{5����}ۻ_GNUfWBd̒_ex�9z���9��Ͱ�	#���=G鸸��d�&I�|!��4���-��|q�H��G:=Q�4):�} ̠i� Y��n4!�x�K#��Q�.��y�ꬥOX�ޏÃ#F
 �o�x�̹���mpKn����5�ۥϛǛ���%�Wow���>�Mo[�#!������`�Qr������s����CD	Pl$HA���Y��]Z�,�T��&�R^'�ZD�h	�&%@�)�`�����?��I ��O�,�,DBHsz�.O��O�_w����2d�$���Q��%�G�K��L>�x��-�}�ǽ��}g&I!���(Mdi�V�0�*h�9�Q^7�"+�&=�I�	˱ɑ�O�8R#��/Jϼ�?H�1泉'��Ϝ���(��3�4s��O}�劣��2a����1X�"���$P�l�M6Nf��7{b��a��hN|�AϏIb(C���(����Ι �-$̄2���O�!��A��P��g8�x>����eW�{,�9� �� ��JX���B4j#���ұfNq�!�rp�	,E�r��,�0(�#���~�#��s��ջ9�� "kW�
8Gh^]���F�h2ς<~��#i���*'��}P��ߠ)A��a�3A/ ��c��{ܔ�݃j��͋
I՝�����6�v�ԕ]O%^��z�9�*�j��ena��ȟx�@�DAx��-���I a��OB�(�lQD�E��B!�IG��SMͱ�%J�BB��$��|��|U���p� �'�8e��������,��&I�ʴ榑�Y��0��`��~��_de�{�$,<�h嚄Yg0��H�d�y>7�wR؁��N(�ܱ	!�<9�YrƕI��pI��QӠ|X���$�sl�$�8���Gi���wF<D�cЙQr}c�1ʚA��G��7۟<(�Q��@������
B�;a��1���q�f/��r*�>(��3�xq}'�9�E����J�3&���K�x��["�;p�<l���M��|N_��O�0�4�!���(�&����X9�?<�7w�:�� �b����������A�.~{�a�E9c�uM�x��lz�f��b��9�}{b���F����>�yF�Ro9Zu�\�q��m=���j�%�q�lEV��I].j�rwn�f]Ubgwe摘)��6>-�K�|O>�S��.=z뻴r9j%��.O����$�)x��k�2d	
J���T͖q�o|i���,�=c�1S�lϦ#nn�k��%� ��1ʤ���B Dhx�ﷻ������$��#�N\��K (�!�s���|ntU;��D9��}�V�G���	8�9x��#������+v��a�"!$q޲-���`���۩]��g1��#�	��L"G� �H�i%����z�zpˇ��k"�$9�2�.X�T���k�O�q�.P��>�N$�r�$} ���	��٤�ލJ����I2HAŹ�9�9S@�2�	"�4�9�a�n���Ssg!2S���;Y�g�!B��m�Y�CE��[�Or�6�{&��կ��H[  ȑ�:*�B������r�|}2��Q�WWt������[�6�a|8@�hm�:�K�cR���ѮC+L�:.�Uq^�w��o��2�U��D@��ąfK�P���b;�GVF�qz��^l2�d$C>�K���&q�z��\�4����|I �i$�X(�O��D���Ey��:vr��S�$�&-� ��	9��-���Q^4��,̭�I'�5�$�	&��� �Β�NZi4��s՟�}��̻Ϲd!�>�ꏤ�NVx�r�p�a7��YOE�$�0xMe�Y�+�Ah�sH=c�#`� ��P�Y��"b��!!��Y�W��(.J"4�Ds�>���_>���	I*�K!�,����0��k�[�1�~�}��|˭���4����|s9x���9���1ͦZ^wɄ�.1��D$� ������ϙ�����?W]ߡd�Li��"Gψ%?�$��X��W������^�I�&�>t��9�,�c
����"DDi$��wD�1%���5(�j��� ����3{�~viӿ��/�xߊ�F�� ����x�4p`�> �)��[�#̨j�vT��:���vf��$�(�e�wf��{5�#f�n��-e��6�V��r.�7G�����<}�<�Z�0RZ�IlL����G�(��	14���-U:V��;�h ��h	T� 	D �#j5
6	e=�
A�0G��ڹ�Ry����`��ş(#�ls����w:&U��	3iA� �$�>$��X��bf�ŕ��F���볘c�6�Q搡�A�'�r�r�4�>ٿE��ʻ��f�I&`q	������c��+��1�s��W��*��`)02m�%�9i���,Eᨻ�6g�=�y�	$�0	$͆H�<d�I��ϋ(C���ƛG3gė��坏q5��]�A�K9D���%� ��9���Y2���C1�N�q��(D�>8��/�:\��aK�w~a�$`�aGA�zJ<��iV�G�c4E���w}����xA� �M-��NZi(xxh��+�\k�@��~5��ǐҾA�<��.e'�t��Ʀ�~�m8�K�3��T���}��g�>A�^��x���Z��542�u]�S��ىs��ݚ$�-df��5�%!��)����� 4��
a�(�A�� @�m�=Dyς!��j��(�	�
)�O� �"�@��4�I-�K$��$�IC�ܨ_�$�����B6WU]X�f�����#��Ae�^�Ћ  M�,��s�S8P�׈%?Ig9b"q�4��2��};�뻹�b�e�I��X�a���Q���?g�J��W��C��Yą���ɶ9�D�� �<�]��,s�p� � P}c�#��8Ɠ����'u�ۚ���5�Aė�Y�.����1s�������U\�68�'�94��<A�C��0�`��Q2F't���M �Ǥ�#���8�ۨ���Uq�Y�G��G�P�a:����On���/�n���g4��9B.	�4��r�;i����/�|K��K�f[�v�����|�X�h�_����u�ݽm�{���yt��l/��������8E�"a���U��,����nv4���Y�u�x7�1_�u�c`�Z���j�����Ftһ}J_6�<���W��;i�;C/^M�z�%WF_�E�c��<6���`QȞ�s���v�-o�jǆ\hf?_�z�����{V�\��=��5��5J�� ����hm�iD}K�_�A��:����s/���yO#J���bze\>�-�}K*�պ.�x����3!�v�<���Y��ۯ{]��J�u=��v#�W&i[��_lB��X:�&�YqUG7�*_z�qmcZ�c�����_�v�i����������^\л�rG
x��h�	t̞��-�>��ǋ9l'�����8%�����[�}�=�ܼ��QE<�#�L�T5�bm5Y݆�Ρ�ɬ?uu��������(,�6V����f_Q���{ۇ�y�_ww�^����ua_���G#祥�Xã3�)V�GZ�kZzӉWsn����;RL�hC���[X�r��U�G��r��GMc��m�݂�8&�����BiU�l��!$w�����9�/<�á�>��=��ѻ����1�H�O�\I$�P�� �$�ꭱh!��Ђ`���wp�6�������r�˒�)$�m���$�^�����$�����Yd�I/r�,�I$�I/m���y痄�	���F� �$�D�5��������A�c��I$�a8��˔d����O]�QD�����b�i0�NۮACk5�cr3S,�=����u�5W+�B����R �Ԭ�lWV��}�J��'z�E�"�V�u1��o���y��P��-���U(eml�.���ܼ�l�4�0̱�Ou�׍Y� �ŤS8ޛ�<�ռ)��ߍ��OK��姑g5�]��n;��jGr�
��!�
ff$7[|,�)�k^\�e�Mۮ.��S���c�N4�QgG6e�fS�f��HU!	�bUt�wS�)���%v-^�MI�z:��Uڐd�`N�ѣO�-�S��w�#U*�]��%r�YEUХe�f&s,�w+�gI�tK#6���j�{t� ��{��M�����:2���!��y����z�6{qv���۬�7Mpn��V�<�����g.]luѸ�9gH}(����k�G�]]��'7r���)��ե�۵�mYqG�m�������S&�GN��9�s��"�o����YK7u��gQ����˾�a��񫺻���+ѳ�H�r9�)%wKp��X!�m����%19�F���W�o�X�.�)=�J�OC*	�М��L���y�&}̲��v̨�N�)k�`(���{A����)E�+:��/&+���"�7���v�r��Ï���<6���7k�y.�q�J�rg���9L�jN��ʨ��5*aBv.ݤV�߬8����.,�,t�oQ�˱*�n��S�mp'7��D��4��4��8�0[nu�
�2�;�\q�2[��m��ٻl�[�C
�4�ˡO-�7Tj��tΜ�j�[��ƴ�ӯ���d]w�$�b��"^zE��Cqle�v�[��J��`HŘ,֝q�6v�ѣƯ's���B\n�;#�y�z�׷�m���nW�^��,w��-3A��n���

�B��:r�J�'H�3GD<�IuN��S�]�uhQ�Y�m/VB[}xh�Fw���=<F��*�N&��{�W+/2�m��dO%�4�+`�i��^���%3VV6���v3#э#~�擾��d;Y���"�iY�E���;vցoY.j�Bhe
OUN=�	�F�mo��R��r>���@�x�N+��gH����74=vI��(fʥʅ�w1��)�)�ttꫡC�1�8Y�� �����8���,m�P��@nm�Ά�䀪Ԑ�ph�yml��ǖ-ʦKuxVQ��$<�1F�i��ʠZ^,�¨�q���&▰��%�A��A�䅐�F$MH��PTn�,#G�(�Ez@��5w�w��-�"0�D_�˖q�<Y'�m>Ľ���C8�%��|U���p�1'>�u���U��s�0���NZi�ab� ᰫ>��i��(�)YhE�&���#��o�0<E���ȑ��K>r�D$�qYe��[��k�י���2.M""��!ܣ&	�p��{�������ݤ("H0�>FpUm�p7�y��ȩ��$��8������ǌi(A��JW����|[i�ĝ�Y�]9A�&sM�½]����w|;�R96��4��daƛF}{��/������[,�X��ď3��O�ͭb�����":��W�P�{���<�v[�������Q��RXwlM3U�T����E�=�݇yw��'��(�[{][xLݭ�#�6}���T'z�����Bг�z՟�H�� �y�%"*�$�Q�N��4��-�!�0aZa�Re�A��M��5*	L& $Y�LRTd���bf[�qQ����&�s��,E�	q�2���9���q�20���M�q�/�,�o ���v�h���dG�* ��Rv�������E�w{������'X��˖q�4�B�`���$��zO��4�<c�[��Zi�!�<q�1��o�}^o#%9��s�,��$a��9����Wf��˻����x��� ���|�	G��_ޙ�w��Y�X������\��J6Nf������k��||I�0H�A�Ő�}�u�>w�]��-#�G��PA�p�-dw����MsqS(�^�C	1���{F[��H��(��wՉ��~>��Ä��|cY�;qV�N_> �4 �1B	-�S��/j-��
�R������;�λ��E�v��OX�z�^�po*g�Z��:f��ϡ&�J��q���[-*p�BI�B��rQ
�4����	�D�OlNjYH���Q�P�dN_�1?�q� N^L��a�4� v�o�j�ʔ��9-˺ DQ!"n�Î}'�9�w���^�ݿ�brh��Z�oAǍ��9i��o�����Uy���d�B.	q�=F�T�����f>����#�5�q�P�+�Y�z�5�9���^c��>�\���N�x��(D�I(�Ow?l�#�(��^�\��l�9�����g]�4�9�U���p�8�O�h/�����q�1�ɜr4��$|A�d[�����~�o�O���>�I�#�k ���Y�G�I,�2����.����c�3�$}}�>'ٝ��/&/���'^@\�/�Z��<�;*��]738p�C�b�lA2�^n^��B�Ke��S��3w�۵&��ܨq]pAMՕ9[�V��f`�Fpt6��k�]��dYN�"�AaJ����`�
1��!+�(6�/�պ.�6F*h�n�״,�$#q�D)!��]�4�:d�B6U�;@V�I�଄�[!Ma%'Ly�܂F���᠎�H��>�˒aA��ݞ|r"I�D>Y$;�l�#�Aǋ ,N&F�?wй��;��o#��PAX�$A�O'4c~F�ѯ�S�H��E�1���i&�c�Ĝf��EL`�� Dx��6AÎzO�r�9\i0��ś򪈏��8;h�q�^�-4��zK8�&�}���̮a��j(��%`�Ń�#���w��3��	��BE�%��X��%� Ø>�g<�1/�S���(.J"�$��f��=�q<.����ßs!�,��}��%r�r'~u���>�%��/�wz����^vf�X;�u`�4�]:���QGŉ��ku꠫����W�t[�}S�
�6"7ƍ���姵��E�6���h�K�1�[�ܛ������D�*D��uj�+��Pǌ�Ҹo05��}@������
("�A�v���'�|�x��a���'ă �!R���m{e�Q�T��$L�J�w�B(Yo"B����{�>!u�������u��;2���p�>�xp�> �O4��M#�4�>��Bw���9��� ����p善Y�}g�}ӕU~f�3�||<���J$~>$���Yg�ww�3u�z�C�I�YpRm( ��"DD4�9����������o#�$} Ë �3���6�G0_�#��;泲Ђ��H�ğ'2� �5�&���4]��g���cIBo�0�|���"8bl�4�>i|&yR8�ɖ9T��8��9���$S3l�9Gt��r�H9Ǥ�#Y��-�)ml]��4�N9�̪RVx�r�8�8�h���S�i5�7Нyu��@��p��/�WP�·�!�-ڇ-�pa���,����Gi�0f�8p�?�
ڻ��x�`ʾK���^�ޤ9]ӝ*t��գz��oEF`�Gr�4�yUz$l�f^ڲF�a@��1Q5(�
Ds�ڼad�CB��*j���u�7ڊCd)���2�sj�ZL�u)(�Ԉ�úID�A-�EzҁL��m�S#�@�� �$�E4�`C���w��b>���ŉ��%��`�s��2��#��;q'��"8��N�9S��8{oiM�U�����
�;�x�J5�-�ҭ4��+�7�ww�1�3�b�eIe���&��<Y��l��(�����C��D\��܊�	,��7�K�'UQX�e�J$�$�X����q�5s�>o{�����57�%����!ܣ9�����LL>�Љ8��8�A�Ѩ�.
��GoΥDc4�_�	"�� slrIv�Ƙ�sQ=���ݯoq�B	n �J�,�T@�<Q!w�ط�G忷�2�o�g�5�m��g��zl�Y��*��C�D���23v�����l�� 4|X�(!����I�O:�L�Nꨳ�վI̽|�7&�y�e�"�T���t��r�L+K��[~A��5ًj�$��A�Wf�Dȣ�e Lm�>F�2<����a��	&*H�N�,��d�aȲ�(�l�5
1�)����Ƴ q��n哕[�`��#��z�]'����&�_9Rm�U'+cP�태4��g�ǈ�f�&M�r�H9�Ib(G�������"�M*�3~R_ØX9BM�8�/3/��ݞ�����a��Q�r�d�xr���N�i�{���r�ʢg�A�|"Fq'�7*Y|id���̩&g c�:�q�.J1�-��V�G��R��+����;*�3�f�� �ǚ��&�Ϗm��x0���=g鸸�5Ԩ4�ȯ�,$��AǇ������d����r���a'`�xIa'�=e��d�G���d��3��&L""�$�r��dZ9�L���
�����Rt|_�Y�Q1=��Q@�Y�S�u�UP��0���y2�`�U׌��f�+y��G;��،o�b �A8Ajt��MS������+�׽΋}�O�`�]�ۼn�W�D�����������Yjn1Qլ���tTcUP��`H�z'Lz�W�����f"�E�=:��D�N׉�"�	����I�;v���������6�#�*�6�9����A_0�gae@������X�������13�0�k$�L�,�˪ DQ!"gգ�p�i�=�Ӿ��O 	c������8;`�i�p�Q��l+_3W|�AϏIb(G���G�����xWL�E�\9���k ��H�W��A��ׅv�Z�+�f0C��1� �r�9T���ArP�`����ݿ��̭`a�x(���9R�sƖ@P�����$LLX�,� �0�.ӓ_MGI����ի��|�f6���9㏰��FI�C�U���|#˪��|����)*y�����~�/m�drv��ZG˺����I�2��42�,A�Kw�߻y��	X��T�bUQ�㼷�V����V�!��U�^�*��4Z�9�B�y����~�W۷�!V�rD�U^����K^��z��x��B��\[S��$0��BbeL��ύS��f�.T�T�Gu)���*'��!��K�j���fU�q���|;n6��x6�ۤ9b M�xy,�Q�c�G������}f�X����x���)6�l��$oΥt�0�h��Yd��Q�L���<Y��+������3<��&D�IT|����z�	#�����Ϣ��5ل@����g1���i&��վ�q�g �Q�{�@�>(��3��qϤ��5���=[�Tfd�}���dj�r ��M'a�S~��*���(���(E�D�|�:�IZ9�����S���F33�6�I�P�z�	g�Ѧr�3��y�����-� ��>r�v�����~�=��||��ϟ^�+��q�#>�<�m���Z���5�@��)i�ɾ���F�S	�[&1[�
�UY�X�88hѣF�a��Aˣ5le������S���5�k�U? �΂W(���R�h��F�Ҥ��LrT�uV\��ܙ��q�C<���V\!�׉ey�� �M�"	����EQ���$^��6׀�4��26��(B��"ϰ�C>GG��}�Bb�m[)^�<�圫սΠ�ۢ������d���`�ß�T��K (M�!l���=�a�T��io�����I���	8�Ax��������-7�8��,,D@��{�YnUiע.�;u+���Ꮓ���4�ic��d#���ns竾ެ-��!�!�QYpRozK��Q>�☱��aC�B(�&D�>8�K8�s�i9��R˻�*E����}c���I� ����{�OK�*�~����4� v�$�r�s��+�K��K�Y!"g���'�9T��A�fV�����5���,���M 枒�Lgq�LJ��M�A~ݗW㮩VܼyL��v�U�J�:ԩ�s�fC��\��(��қ��QϮ��y����\�_%���(#ផk�5	�5W{��Ѩdߊ�fA��s�YJә�Y���,m|r�]��y6�5�2g��`�m��B���
X���g}�������������jӏA}�Ic�N��*ﲇs�k�ln��r���������ܽ�����1�8`W���}����NIZ�8�v=+���#�����Z�\u�g���/��jy����ь	w��s4`3`�3.�(��T}���VnW�&N�z+�}A�4'�A\��7��,�r��ߐ�:����e���VyR�[꽞>���s�ڽQva����ͽhl��{R���<���==�q���<�cJ'2y�YM�T�?t����X|M*�h��#��'���P�<G-����+���K��w}]Y����^E��M9[��_�5����+�=��3r�#r���!�U�s��Fwz�|��h]}>(ؒ�)\��/���2G]QKbö9����g'��L����5I�qN����F �꺣��Y
�`-^�p��w�1��˜���M�bӝ[0#u0Z+-�Yy�-k�G���r�<�v]����� ��l�I'�g�����}��h�� �uӜ�����s�� c}�'w- �fUVd̒H ��AI$�\�m��$��m�I$�[m�}�ޮ���I�$���1//,�I%�ߵ��m��-��d���,�I$�\��d��.��m�I$�L�T�^NAe��I$�]��n�L�$G�k�24 u��E�d�IF���ڦ�X��	qT�C�-�p^���������qM���v����nn^�t�%cr�$�����8�l��;��]�Z��^h���0����uN�� ��.���/o�F�����;Swhe�r�J�<\Y�2�ڥ4�ལh��RV�������F�{5�:��� �yvN�f��^�sq>�,�d|��A����h�aP����B��uZG8�,S��w7ݾ{���)[±ե]IL+j��E>묧�սd���}�f��[�.S���nR�47&뫢����\HI�	�_p�G)�v��>:����M��2�:�k0�]m�e-��!�VU;���yqy{���Λ��':�umJNl�Ut�:��k�|��#�������Q��v���j�oe�������X[����K}�� ����{W]LMu���޹WU	)�n^q+��(;���T��
�vV�w7�t�環�J���=���댮����b��7��ٕWS.�tv>z�u�F�Ul���^5�RH�E�7w)l�0�xD�)p��<�D��xգ���e:V%hE�rV@�Xے�.�aouS�w(i%Z�(3�&{s==�0�\�H��:0�B[Je�W��K�}��#9�#��>un�J늓�&�)�W1�j�)��ï��u�-ƣ�D��[��WU�]�N��F�'I� �b����y�U*>����6R�e�D��"d1/2�Zf�o�v�YQY���n�n�4��D1�B��,5)��gL�l.��	�uh�����K_aw�)���R8������\� �ӧ��c���.^.�D[2F����j߲ҏeKs͊ު�(q�&����I�s[A�Һ��V�7=Q7��4R �s�z�0ѣ�+���|l�|F5�gJ$9�v���Ӳ��z���)�l�����ǰ�b,��KUb'����Rݕ�6�,��9�
T������#)��̞���s�x�"0��=��*������ͅ��u�Vs+��C:�h����B����N��evb��9��CĞ�$]���@�v![���5�K,�l��*3*0R�U��B�8ٲ��w$ ��{(i�g�%�mh�028h�@��A�S3y���	����T9���YRnj��}�CU}�]��U����s�X٭m��ieWh�{��@���x@���N��܍L�w][��9� $�?"��D3��>�g���/2(��	HH�E�x�uy����p/b˘kĂ!�U���IoiNK��0�/�r"�����<XAB?0}��{�e=7��qeBE�%�����& À��u#��ck�|��%� �$���p3����v���}kc���Yd�	�#IF�v���O��������3�($� �,��K��&��4�fM�����H��H�	;��ܪs��H,��gy׽q]wz�	�4���|�	������#��^/�⻻�xᏥ'��$��&Ib$DzM�9��V�1�&f~dl�"�>,���&Fx��f~��ÝU��9��9�8II'� �,rIv���D;��ޗ�N��V����I�ǅW��x�2�׺poS8|����>?Q�U�6!���{FI�Gަ80���;�3M��l0ŏ�h!�����%�\�1j�r���O^&*�]vbzc�s}o*hNb��m%���̩M撫5n�I `h)q��x>L�!~��,��!�^�R�WC&z��&�^#iy�a�$��B)��Or�,#�/A9qwfc�]�_����O���O���Ӕi��N��/�&U=y� �3���2M�ʤ�q�5sJ��|�T��L�<aę� ��|t�"�pW׿J�z����|%� �q�JJFP�a�M6�>$�}��9fDօ"����A���`� ���!�|aœ.�-��,=%� �$����i+���oMU{�0�$(M�!I�<���V�O0^�����+�����im%�r�H�mX�3g�;f��U��0��d[�Nqa$"�5�����]L��9����	���;,C�Hs	4�äGjlz�������ߗ�  �|썥�5Z��#������Gm]	���W����'Pj�|=�}�4nKP�e���:�8Zme�w+r���`�]r�d�:WJ
������u��6;eɯ����-�;[7��S�Ԍu*�ܶQM�r�5v\��U�AV/f/$]!�ӗ5B�'f������3\�&�AIb$Dl�I��'k��T���H,�,L�dx�M�Q�9uG���K�X�P�$t�A�X��1��o���N�ٹUy�� �K��<��"Hp=�����U_xM�)s�}c�I����8;`���gK��ux��H9��X��K�A�ѳ���IuU=�gO�L�s(C���OBE��i�µV��웿��Y� �Eȉ��5�)�M9�ܟ}�j��o�B#�0��}��,�4�dsi�-Z`�k�B$���]�*�,$�������~��Ɵ#��B��O�:�=�,�("�ɫ�A'J o&}�"�	G[��^�����nu�(�0�#��6hK�9b]��/���֧Sb�4�r�ýu//��zR<�e$o�a��7r��^'u��#��3j�e�m�m�f�0Ez�أK.t@��̜}Y��(���!��B���b�p�T\�ԗ�p�>o�8h,�x�d���#8c
��������	�
1ʫ ���o��GNg�f��ls�{8���	!�$���ይ��5�
���&���DH��>�F9$� �Nf����n�}�}�zx�&q2$�̣�a�]P9���^z>r*T��<�qD9�9$�|q�Kpt�{���\W�[i�ĝ�Y�]Q ��BD�壎}'1�G�����˻��NU�A�C��|I��#���Kڨ��G15��Ib(G�K�A��j�����>&]�O�(��i��z���PK9�gO_}_/��b�.����ZV{�J��4�S7���\4^R2F�G��F�Gf_:��֭zj�~�׏�1���!��v[���0��V��R\��y�q<��լoh�e��TjG�j�`�czk@�']7�a��I΁�̹y.�"��)��d4��4hqULqdA�cM�Rpw�4��c��A9�-S�%������E�w{�9����,F��K!�4�
�s���3
zD#O�v����I����i��qo�z.�y)̑��,�0�� H�	7�s�qg}����ww⽤	�&���y2�"G8�>�'x�x����������PA�p�q��<u�M9���|9$"���M ���,G3I=u�?}��v�����h�1˪ ��G�Lf��1>� ���]�Ìi,@�$�b��2��{9-˺ DQ!"g���>��y�ظl���W�p��:��hM0�6;�$Ҙ�/
/R��o����!��}�5J�I�q�h[��(���m���0��hD�}'��b��-���5c�5��W4��e�J���矠7�+��h���UZ��M�Jp����xA�����=m������Lٺ�^"c��Tƍ�����S�PW�}ӋY��ͺ��cZ�oi'�70��I��]�o��z���3�<GB.	q�<�6�IZ9���1�o���0Mga�$_ʠ�s�=c��Iͧ�o�����B4r� �QN�x��,Aq�7Y&��~��G�P��ʖC�,��ǠB0��s7�Va�d�x����XI48AA�xr�����q�<���8�4�� H��N�,�*�������l���ｰx�|"�\�<��ȑ��H;?0g�����SW�g��$9d�A�,����k�w���L<�ÒB(�$��<Y��L�=�}�V.O�;�]���i쁟H����O�^��K	8Z�_�E����������z=*�n�P*鞼���h�U�([,w��5������w.��l�+ꊮ�kʧX�\����HD�F�nV���R�k9Ut���A]���$I��H�Z�t0�j�̄Q(��T���h�%[:��n�h�_�����r��H�OA�Ϳ#���ڊ��8�ݨ��4� v�H$݂�s�$~���D"����B�A袩9\i0?i�f���!7���I'^�&�sOIg0a<N�v�U����{��QE�)+��P��w��DG�����㋡"�T�i�p�6DH���v����~��#q;ae�B#�N(��f,�n��wwoƜy!�,�
@�a&��]�9�����}�&�L=�Y�'���p��ʑ��l����}
�˞0>�#H$���r��,$r�/W�V����{��y�7�Dz\b�V\cߡd�E��<ۢh��e.KiIk�����z-Ҥ����0���2�;�2)n`j�v�W�DDԾ���r���̩:��(��G`�uI��5<�yB�^Լ�my�4�#�� EAu�xBW�TY�t�f���>�(\{o�$�������X�x(WnX�ﰳ��ݝ���}I#�$��e�6�zK"#d��#�����&bp����H0��,L�da��Q�_�#��xOGx��r��H�<Qe�I.��7�v3>ϑc��P���$�Af9UD�N ��(�9�EL��*G�2�*���cP�}���L��cX�a}��A�=%���v�nq��*�^�#H�̪PU�x�r�8�$�h᠓�4�ދ��#��[��z�(DzD@�A�s�U��$B�cq'��ğp���)U>�|z'>%��U�b���F�d"�s��dm�Ѣ�J�C�Z�+�f�5�<��ĚHI�RKZ�[�q�kq�7u|E���'{&���b��2����v�{|��3�|u"���V�̵�+�I��2���eJ�ЇMk!�5&)L��Y*�`�\O���Sd�q�$��
�O��]�*��DO6Q����/1�3���DE�A~NT��i�d��8g���Q1�s���"H0���r�,$r�@���Oꓪ��h��ǃpr$q�8��9bC�I�����s�?���}� B(���PArX�'�$�Q�sy>���C��� �8��8�i&Ѩ�������b>>�E��@�����1��j'�������"t��Q�pY�*��x�C���/~�ڢ��F��|8�I�9T��<A�C��i���y�x�Ƴ�'~ ��a�X���(r���y����Ī���=�ٍ����o���|�-�������2X�F���J�K��	>,x1a�_����X�°`�4h��4h�{m���ƞ��Y)c��t�[v�7p�u�6n�u
�Q�m�F�e�T��XX':��z�>G���R���	���wg.NL�;�^����6�lwg<�!�<$��J�S��i��Pa�A(�a`$o�|x0�~~�8tm�Ñ��z�(Dd���A�*���Q����}ʓ�3�\�Aatqd#�r(1�ûs�D�������Cpr.ӕ^,�D3Y��ۻ?GeUfp|\�}�� �NT��|x�0�� H����q�v�eG�>r��	�&��8q���G�d����r�~0��r�<$�0��Ek�ux�#�u���d�".O�$�Q�I&�xㆨ�u���>��_}�8�3���mF�U�m�a�aex�A_y�ǎ8��;w����t�翍�f���f���6͇��������8��l6��g�Vm�͇}�cfۮs��0ߖ z�����fٰ?��M�l?�fٰ?���������m���o_��?��ߧ�����6�S1�a[mLeՂ�b�[b��kdkK������%���mY�fl��aXPV�V
aXV,+
a&Յle��h&,!m���� ���XH%���¶ڰ��,!6�L[XZ�ɵ�XYa ���ad�BɖB,E�B�$-b�E��[X�2hE��!mmbe�,X�5�����4�lX�!al�6�1bŶ!6�̱3!c,Y�e�����,жB2��be��,�b�Ѕ��X��-bЉ�ŬZıBЋ�&$,�kb[E�b,E�!��2,D&��-aX��š�[��,V%�Г&�k�X�(V�LK	bе��D$+�bLZ�X��BhYb�b!bb�e�$,B��,[Bŉ�L��hAb6�a5�2�e�L�k�l�f�l��2,[!f���ڶ��F�����QYZ�eUKRҤ��IZ�*R��J��Օ�+(���Ej�b��5aX%Y�X�aM��S+jĶVj
elVV)XP���m[SVڱ[V�m���lSVjڙ�efP����cV5���mX���mY����m�cSmCH�a[j�LQ�e52����*J�թUJ�F����*�+5mFVVVZ*��Z��jښ��VV���m(VSV���*Ԣ��)TV�"�UF���R��JY*R�Q�)E�����j5M�j͕�[m[f��6��+m&�)Z�U(���ML�L�j�IESVIJ�cQ���V�0�$(�[2�Cj��aXE�M��XZ�XZ�-��������mb�kh-��m2bb	���m��-����ma	���m1lXFh-���fXL�am�al�mam�,AXB	a,(+,XZ��V�e³-�5���m��&�9�XM[jٶ+[kb3XY���5�����ڳm�XV��%����� ��k-��AcX@�����X[m�&e��M��5��X��b ��X��XMam����ѵ��A��mmam,&��m�X[,&���&&����E���XH%���kXK�����h-�,���Ya#XF���Űi��6�����l��6�XX����	��kXP[XVڰ�
a-� PS
V��ژ�0H�X+
X+ad�XKXZ�ɵ�al��X[,-6����KX��Ka-����ń,!6�XAaaaaf�CLCXLkafh-�[i������Y�,&m��͚�ى�42�am�XX�Ma6��ab�Y,-�&��6��,-���ml������a��1��,��Ѭ-a4��[k��ɋXZ�H+,,����XZ°H+
��4XE����kmk��Ae�k5����e��kma�5��L[k2��XX��6��f��e��afXFAl��ɋe�����a�K	akmh-aLZ�[i�+
���Z������XPVڰ���¶ְ��XMa[kAL"¶�Ae��i�Amkk�Am���a6X[k ���L[XDamaam���aذ�k	��A���1l��kmfXF�X[cAm��Ѱ��b�m�3A�maX[cXC[l[k6X[d,&XZ�M1-ak[hAkXYa-�Ak	�Ŭ-6��XZ� ��VXK	����%����(�Z�[i��ae��֘�0���m�V���4,-���&XZ���XPV�?��~�]�f�������ٶl�?~?��}�[6́����l�6m��L�f�����3?�6f6�Ǯ�o_{�קn�m���ٶl�ߟ���0��0���3���?������[6́ש��������m��9��f����?���PVI��E@�� �w�@�����d������ �`J�v�������<�@]�ހ�)JQW�7�P
�ܸu����9�#0 �]jec��iJ��r�/ J  M T 4   1�*J��Fb1 �`F�  	�`E<ڃU$�4 �  @ 	5#@�J � @   �"��*~@� C�z����mFÛ U� �@EK( jMb�v*��[���ψ�?Xe�H� E��!R�"*^;y���vhTI2DQH�m���=,5w���]h&tTٜ�uJ�o���`CI���R����R/ֽ�2F]0�H�L�e�K��C�W��.�ɋ�jl2��MMۑ�$<�z�ĭ��8o!өf
��z��	��0�,Za/���!2����:�.�+s�r��ɥ:;SQ��_j�rf[�V\�R�՗٪DR��M͹��Y11Ff��Z�d�+)n����hHS�!�S;i��@����%c(�L�����Em�xh����P�o�vq�Yu�f�4�ކ�8��ݸ�ps�"k�wJ��<����e�Y���.�8����16̹ۉ�.D���Da�A��E��<�l^��e�?LJbES�bYJ�o$as&k0�eI�$�nb��̹��2�f&́��r�
K7x��P�ɴ!Q6M��NN;W�흌����Y�wUEnT�˸���TT�"T;���fԆ$�Ĳ�}��f3��v������d:U�F:��U�G1��0�%w�h��r�T�wn��b��s�L�N)���8pM�T
�4� e8�R&,�&�7j���3#Y9j��*zt�O#�9KE˔$0拔�<�=��{����=��F|^V�s��d 	���2�� @   UP             ���          ��   �`                  ��              �`3HW��w[h �]�ٻr���`��y�W���u�"��)�9�S��N�b�Ewruڒ���kA��j�+�N��6��ՙ6{j����I�&�d�e��KS�v�-F�#E������&��	���v��1S��Q��cT����ྼ��6Pڽfj
`��"nTQ��m�b��Ob��dMi	yJ�MFϜuoK(�t��RC�+���\�Ԫ���I�o
�^ڝ:/�%t�ڴ�U��s�x�ܼ�� 8*�GIw+*wM)4�4��t�J� �θo�7���%����]ϛLwwv��������\W��QU�r��<�+�no���iw+%��,wb�v��U�U	m&���u�J��.����oD���ƕpT$UR� 
�R��/c��HDøQ�^�{Nbz��sZĂ�n�aR���{�,M�0�����*&.n�E\�c��m��� V]��beV�i�X��	��R�YN^����%�u��0�u��K��*E���u�Kٙ��B�C���  "!�� besa��LLm�ʫ��j=�$zȚR�b��3r/+��Lv�d��\J��qKs�N�r9{���K�Md�gwT�\�Q)F��bf�]�n/��՝N\�OXŮ�S�c(M�U;�w��K����i�6aW��qI��������6��'!I�[�\M7r^ʻ��m�$��|����j�ڑS�e>�q�q�Gwл�Ț:\]��z�ʤ��	S�%��nE����K2H�E��'T����Ȁ�^"01Oh�N���H���q%7SMl+����6l�4|nmnQ�iIw�vYY<�uFy"2�JQ8�է7��<	R�"���d��T�!P�����2�I�ab�����
��d��+K��8�M��:z-oZ35.���hy��{ǶD�O2g-���oڢa�5{�V2]Sl��3�N��0��Ur�^%t�-���Ғ~)E�S��ɨ��'���)�..�&�KN�y�]o������={�lSX�r+&r�mwj�]RE�O`��JB�m$DLDYέE��{����{���� �U�L���+��#V��[��9�h�UEϝC��B�H�4B���4r��ku]�7Ou���-�$6�b�(��AiDX*�����/x���P<@�i>�ܿS�Ș~{p����8�n�r�w���*�2�V�A��m�J�GY��+H��1��6U�͟]V�6A�p�,�J��yrd-��T�Vws���4�Do7�_S�b��*�o�������y��۳L���ہu�ѣ��'�*�]�o��/c���u݆dm"-�g	��a�fn^�{ى��^>T{D�h����Z .A���D)�i��=|���d0�kR�&4 -�tJ��4��DE�R��v/9�Ax;Zl�`>1l�ɘ1�e4�r��"3G5�/�j���(�������ڢG1'p�\ �{��/��gΦ���.	p�|��D��Q5�FZa����:�o(�0jUC��5���g{>Mp���� ���l �5���6�n�up��|���D��WNY(�8�k6��SQY�=���e�ln�����)RR,���Jp�0STR�)b��UGJ��i��ybZ��hU7�z��:1���p���QG��΋����_Q�nj��k]��"a q mc
B����-�0����`��Q4�&K�G+j�!8�@ ��Cl�4�7k���o��ƾ׾+�`0��No�$4�)�L�@0���d�@�	a8�L&����Hi�B$� a�iIa>�`�>���C�e�f��d��'_�����{����U�|����@�

@H w*"&���녗Vō�����)Xq4�~m��6k|�����@�Q�"�QAf�F�m2���n�x2�Z�Y��}T��uE]SIH
�P!�H`*�@IVU4�B�U�Ȋ7j��o�v��-�(o%v�{X�GtN&}�Am&S��e�m��t���I� !<+r� �V��PI�ʡ��w��E2�>�e�RN��铛��y-���ޱ�����ɠ��NNd7wuMKT"8PArn�Ai�Մ:�8�2�%�E-�wV��wRBa���� J#�1R��n�˙νr�B��)��r��C�[6�!�L8�`��m�����CiM������e�%0�/�4���P��۳|؂�Ob�I)4�$aOKa{�6�����7��t��y@�ArH�h�$�����D�-��gW{>�g[� ���J�Z��N���f���źz�C���F�hdQ3l H  *��(*�����q}�׽t�U�o���/4�
���K���ɋ�2�r�N,/ =w@�N�B�Ȥ)���׼c�}���E�+L+Uo5SH�����2��~�mOv�0�ZN%�Y�ѻ,�h�����|�7��!��Y0�9w�C/Y�eʡ��Xe2�4m�6�C	��i�ַ�u�Y�<G�������$QG$��(E�����Ұ㗻�m0�j�KN��)B1��D�i�ۨ�ט�0�"�	���T6�M'P���l4��L��O;^T-�S/RV�(��A��y����r��$$/0��L&٦Ze��a�>�8ɯV�[H)��h.U9&��s��s��q��8�� ot[:����ۗl��⸔��Ro�ċ�I��s=��}�^op�6�N!��C��4����˥�:v�E���3H��N�o���w�[Vi���SIĞr��b,(O2e°���~�������m�0A R �t��u|NT��d2p��,����L�x������f��N���9	�!IA$i���wr�6�"�9�ӄY��a�N��l�B���2�o4C��%�����:�Ru�ݞ�޾,V^Uu*�ݡV��[�m@�>^ȩT�0CS�������w8����U�����J�ގ޻Z|� ���� <��ݲ�^bӮY�����D�����zD������ꐆ�bN��������i"�r�h)E�PbE��V��[���Ʒ��[�)�0�+�e�L�18�9x�S��	N���z�,Ɋ�JIl)̜�=��ݫ�z��Pa�*�D=�h�,��cU�8i�]߰�M�\9`x#�"h�c�:\8��0�Ѳ����	�v�풍F�qg/�=�r�D>����{��,F��ڍY�`���Iˎ�F9%�X�s��v���5k���ވs�'-.���U�!��s<�9R������3��(od[��Y/(.l.�]����f��S��؁S���� B�6�r#��f5��G^Pb�k����)�Z���Ntճl�d�:0�h�u׳pk9
�lz�M���s�N�oGr8�f/9�1Q�hEg��m�VG�0�6$���*����!�+k�3�՝x<��x�34^7Es�o�9���mkg�ǭOV�â|6�      @L�"������Z�C�k2ys�^�ɘW+O0�DP��	�Mm��m�[�7�����v�LE�Ȱ"ÈP�e*e%Us���9񋽯���Y�#�f��M�w^�� ����>?����,̌�E��vp�]x#�j��[���ϻ/��5;��(u� ����*uB�:=chi���Mdi�:0��w4���d�
�Ҭ��znV#�;�9^�A)bV�G3f�J�Np"	�y9"�G���nެ����@kҬ�NT�������iġt�z;��*�oK�0�%N�3��ah)�KH�
H�DoX�����q�����Q�oiX�n�Y��Pu��^��7��(D	�]0�������AEn� ���F��A!��縔�]eu��O�s��������%��:U���l�5[�s9�JQ�G�R��X��%���kh�j�K���ʬ5+=�t��{\z�)F��z�`����{c�^8B(�ά�-�` UQ��  J����-AJ�v+��f%�m�験(�tjo,�=����18��(N�Q�ym*z�H(�i��(�Qr��fox�����oX��Ƶ٨�`Tmqϐ��#�X�OGv��wd`�g���9��;�b<cҒ吰��b+"����S:
V́���6=jg9�yZ7��\e�X�c����d�N�	���r�s�w]g	�5[�Xî1\�ֽ/��N��u�{+qt]^ �h�/�}p������� L@ikzr���S4�_rQ��joiVm�C���#w�t�;ȜY�
"0	��gX���4A|��c���[�]�/77l��ہui
�Q݌Q�`����o}]�&w�nV�a���Xo�#�yԄWтr2�|7=��.��*�ڼ���y��aN�W�A3��U�{��ڛ����fYw�մ����E  �   J��Ji)�sϢ��l:�_Ln��y��]`R��DIR%DUf�y�7��w�k�0���qEb�"
����A�2R��UU*��)��9Oźp��٫,���"=�D�Kǒ�;�H�2��yk��<)��HR)c&2�ӝ�;A�Bڹ�j�P�Ȫ���.�����b��޸1�m&�Zd��Q����u�Ӛݚ�����mF+����F⊈�U�7,�d[��\Y�yfnosR]�n��F���Sވ��諝M��;�	���P�u]ƭ)��`gq�mM��rEp�څ@c���*f�@C�\�'��W
��	ء���yU�,ż	�wl�6�aY���§qq0�	<"<�+�=)򓽾mf��.45"�zȆ^��sR�DGOw���z����]�M@��*ͳhw��3���1`���췚��<P��ve�M`�ɢD�ZW��̋ǝ�C���n�3٢o�+&��щ�&�b{fcK�e�O� ��1�  �%U30���&4����SY�Q(�Q�c�+1i+(����s2�cb72��3U���*�JDX����b1��RR ����Z�y��3�w<�E�y�7�Dy`@�4�/���>*��~���ǰ�s�1��y]������� ɨ�A�4�3kw�1��,���vaa���L "��BsE����蘌�c_w2^(3�و��m�57E�T4����C�Gz���F�7������缔e��������s{�o���%W3�{��+���{��!W!����JQ�s�Ć��5�Y�x�\x���n�Ձ���IR�\5����݈��A��"9g�k��}�5��v��PU)&*��ީ�F�������	Ew�^s�b���8E�|c���f/��^�6�H�QQ�V*
"�F1	(�$�JR�TNS^��S�I����v�����D�)L�y;W����OJ���DE�
*(*�I$!�-T�5#��":�֕�g�	_M�8v�ݵ��Լ�`������ۀ��6�fN�C:�4yڱ뚹wk���뷾�]ѳ=�u<���ʌ�X�wU  �@  	U
RQ*�sP�oo'2����i8���l��*�R��IT�&E(�PF�����f�N�LT�E"��"��	L���
�)99�V��ι��qU�K�)�1��aH

JaBE���a�7�^s�fb�n�q�&=�xu�>{�/�{��y�b��fR�,Sm	EZJ����D�����q�d@ZG#��}�����=���j�m�zd�XU
@PK
��JZ�RQUH��J,�i�;��N��f��6���ҵ�xt@�B��ƫ]ǻ�o�5US-"��`(�Ue,F2�<����~�5w�8����qײ���W���M�U5�9�&�)Q�R�)�b#PV0t��o5z�/��s��a��ӢGw�E�{d�-2�K�@׶A�V(��E�P()33�b�4�/:���-M=剱���+yw�wڮ���a�b �_@���D̫��Վ�#"xr2b�lqh��O��Q�ؽ��Y�9��'��LLQ�T��/��N�h�z�{�-5�/S62ӫA(��S�&��b����Y)E�ɼ�m��¨�R`/D.���\Y�8ʩ٨�8���`f(�<vD}e���L������nN�gle`�Ϋ� �y{�v���f���.�H��W(R�����2�n��U����� UFcl ��A5����2�ˇ�1<:��h�Ww\p�_�^}5C�ܷ���i8�p".}2b�&نe&XTB���������&�%n�����&"����Ol߅����j*3�����8��<�gX�Ϧbv�Xꆅ�\�DP���X�Gs�|v/o���f��WJ�k���������-i6�1�j��cܐ{�G&4���ӄ§��$��8@\�7>G�e��.�Ua��1���֥LwI��p�D�K7N��F�]�5[ǓJ�dM�6`�� �%�
�(���m���zkO0�G�����4ss}�w2:ﳫq�2T#�t��Xg5ۚ�8�q0�|�7��=�+�=\b�^։�ۣ@P |��D	���6� V���Dj�rP '��S�:%�9Y��h������5��i�(�k��bQ��+�Cw�i$�I$�DQJ��E;�Խk�B"�//�p[�,�¨��ƔT(�����H7��̆h�@QW��,�Z���wAE�	�ֽ�jՏ���C�W�:s_��oZ��>-y�KK�E/���dtb�/s��5����_�(d髬� ��h"�z	����8�@�i�����0��?��m^}K��E2�<�r�UŠXn�YR!����]�ၰM�Ԩ�-�e�CM��u�")e�(l�� ��dP��@H ,���@�! �� X�@ *@ 	 �$*�`� �D ��20@P Y@$T�Q$EXEV	@$ �P$Q�@^�@,���@�L1�s��\�-�r=QSQ�7�[f<6��o����t^c!LM,��)�����""�o�q���������ܞa��M	K���1��^�ë7���x(�aγ����w�A�r�p_�a�N* ��y"(��>��!р���B����-�.�D-6�d-�vy	�PT�m��o����pB��s ��.�����hAS�����l����?-���܅��������u�x"�v �������������ç#ٚ��ҹ�]i)�#�����g��8��mSj!cˡ5��`�P����`�u�
�7(���N�ǰ[s"xjQN�z�U���(�LV�q�P��]$�טe��"�(H�<�